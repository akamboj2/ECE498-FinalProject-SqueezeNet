parameter nbits = 256; //note this is actually the precision in bits + 1 (includes zero)
//^note this is only in this file. make sure to change ram file and testbench if you change this value!

module fire(
	input logic reset, Clk, 
	input logic ld_MAC, //these are control signals, currently i'm sending from testbench
	input logic [7:0] in_input[9],
	input logic [7:0] in_weight, //only used for 3x3 conv where all PEs make 1 pixel
	input logic [nbits:0] bias3x3,

	output logic [nbits:0] PE_added,
	logic [nbits:0] out_PE[9]
	//if this module was a part of a large nn there could be signals here indicating where it is, when to run, etc.
);

//logic [7:0] out_activation; //inputRAM and weightRAM output wires, outputRams input wire
logic [nbits:0] out_ram_addrs[9];

//here we should be doing 3*4 = 12
//PE PE1(.in_input(in_ram_out), .in_weight(w_ram_out), .out_activation(out_activation), .ld_MAC(ld_MAC),.*);
PE PE_array[9](
	.in_input(in_input), //9 different inputs for each PE
	.in_weight(in_weight), //single weight broadcasted to all PEs
	.out_activation(out_PE), //9 different outputs for each PE
	.ld_MAC(ld_MAC), //single ld signal broadcasted
	.*
);

assign PE_added = out_PE[0] + out_PE[1] + out_PE[2] + out_PE[3] + out_PE[4] + out_PE[5] 
	+ out_PE[6] + out_PE[7] + out_PE[8] + bias3x3;

endmodule


module PE(
	input [7:0] in_input, in_weight,
	input logic Clk, reset, ld_MAC,
	output [nbits:0] out_activation);
logic [nbits:0] out_MAC, mult_out, add_out;
multiply m({{249'b0},{in_weight}}, {{249'b0},{in_input}}, mult_out);
add a(mult_out, out_MAC, add_out);
register hold_MAC(.data_in(add_out), .data_out(out_MAC), .ld(ld_MAC), .*); //to initialize to zero hit reset
RELU activation(out_MAC, out_activation);
endmodule

module RELU(
	input [nbits:0] in,
	output [nbits:0] out );
assign out = ( in  & (1 << nbits)) ? 0 : in; //if in is negative = 0, else it's just in
endmodule

module add(
	input logic [nbits:0] a, b,
	output logic[nbits:0] result);
assign result = a + b;//(real'(a) + real'(b));
endmodule

module multiply(
	input logic [nbits:0] a,b,
	output logic [nbits:0] result);
assign result = a*b;//(real'(a) * real'(b));
endmodule

module register(
	input logic[nbits:0] data_in,
	input logic ld, reset, Clk,
	output logic[nbits:0] data_out);
always_ff @(posedge Clk)
begin
	if (reset)
		data_out <=0;
	else if(ld==1'b1)
		data_out <= data_in;
	else
		data_out <= data_out;
end
endmodule 