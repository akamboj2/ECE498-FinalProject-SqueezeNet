module tb;

real inputs [2304];
real bias_s [32];
real bias_1x1 [128];
real bias_3x3 [128];
real weight_s [8192];
real weight_1x1 [4096];
real weight_3x3 [36864];
real outputs [2304];


    logic clk, rst;

    always #20 clk = ~clk; //generate clock

    int counter;
    real index;
    logic signed [7:0] val; 

    logic signed  [7:0] PE_inputs [8:0];
    logic signed [7:0] PE_weights [8:0];
    logic signed [7:0] PE_outputs [8:0];
    logic signed [7:0] out_3x3;
    logic signed [7:0] bias3x3;

    logic signed [7:0] output_s [288];
    logic signed [7:0] output_ [1152];
	 logic signed [7:0] output_3x3[1152];

    typedef logic signed [7:0] logic_da [];

    logic_da lookup_input[real];
    logic_da lookup_weight[real];
    logic_da lookup_output[real];

//	logic signed [7:0] lookup_input [real][256];
//	logic signed [7:0] lookup_output [real][256];
//	logic signed [7:0] lookup_weight [real][256];

    fire dut(.reset(rst),
            .Clk(clk),
            .in_input(PE_inputs),
            .ld_MAC(~rst),
            .in_weight(PE_weights),
            .out_PE(PE_outputs),
            .PE_added(out_3x3),
            .bias3x3(bias3x3));

    initial begin
inputs = '{0.125,0.1875,0.3125,0.125,0.125,0.1875,0.3125,0.125,0.125,0.25,0.125,0.0625,0.1875,0.1875,0.1875,0,0,0,0,0,0,0.0625,0.125,0,0,0,0.0625,0.3125,0.25,0.5,0.3125,0.0625,0.375,0.0625,0,0.0625,0,0,0,0.0625,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0.125,0,0.0625,0.4375,0.125,0.125,0,0,0,0,0,0,0,0.0625,0.0625,0,0,0,0,0,0,0,0,0,0,0.125,0.0625,0,0,0,0,0,0,0.4375,0.1875,0.25,0,0,0,0.1875,0,0,0.1875,0.0625,0.125,0,0,0.25,0,0,0,0.4375,0,0.375,0.1875,0.125,0.125,0.3125,0.0625,0.1875,0.375,0.1875,0.25,0,0,0,0,0.3125,0.1875,0,0.25,0.25,0.25,0.4375,0.5,0.375,0.1875,0.1875,0.1875,0,0,0.125,0.0625,0.0625,0.0625,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0.5625,0.125,0.375,0.1875,0.1875,0.25,0.125,0.0625,0.25,0,0,0,0.25,0,0.0625,0.125,0,0.1875,0,0,0,0,0,0,0,0.125,0,0.3125,0.125,0.3125,0.3125,0,0.3125,0.5,0.0625,0.3125,0.125,0.125,0.3125,0,0,0.1875,0.5,0.0625,0.3125,0,0,0,0,0,0,0,0,0,0,0,0,0,0.0625,0,0,0,0,0,0.1875,0.3125,0,0,0,0,0.125,0,0.375,0.1875,0.25,0.1875,0,0.1875,0,0,0,0.125,0,0.0625,0,0.0625,0,0,0,0,0.125,0.1875,0.125,0.125,0.125,0.0625,0,0.0625,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0.0625,0,0,0.0625,0,0.4375,0.4375,0.5,0.5,0.0625,0.25,0,0,0,0,0,0,0,0,0,0.0625,0,0,0.125,0.125,0.0625,0.0625,0.0625,0.1875,0,0,0,0,0,0,0,0.1875,0,0.0625,0.125,0.1875,0.0625,0,0,0,0,0.0625,0,0,0,0,0,0,0,0,0,0,0,0,0.1875,0.1875,0.0625,0.0625,0.0625,0,0,0,0,0.375,0.25,0.875,0.125,0,0.375,0,0,0,0,0,0,0,0,0,0.0625,0.1875,0.25,0.3125,0.3125,0.5,0.125,0.375,0.5,0,0.5,0.4375,0,0,0,0,0,0,0,0.125,0,0,0.3125,0.375,0,0,0.1875,0.375,0.0625,0.0625,0.375,0.5,0.375,0.25,0.1875,0.375,0,0.0625,0.0625,0,0,0.1875,0,0,0,0,0,0,0.3125,0.4375,0.1875,0.1875,0.1875,0.375,0,0,0,0.3125,0.125,0.125,0.0625,0,0,0.125,0.25,0,0.4375,0.5,0.5,0,0.25,0.4375,0,0,0,0.5625,0.125,0,0.0625,0.125,0.125,0.3125,0.375,0.3125,0.375,0.125,0.25,0.1875,0,0.0625,0,0.0625,0,0.1875,0.375,0.125,0.125,0.125,0.1875,0.1875,0.25,0.25,0,0,0,0,0.25,0,0.1875,0.375,0.3125,0.1875,0.25,0.3125,0.0625,0.0625,0.375,0.3125,0,0.1875,0,0,0,0,0,0,0,0.3125,0.125,0,0.125,0.0625,0.0625,0.375,0.25,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0.0625,0,0,0,0,0.125,0,0,0,0.1875,0.3125,0,0,0.1875,0,0,0,0,0.125,0.0625,0.0625,0,0.0625,0.3125,0.125,0.375,0.0625,0.1875,0.3125,0,0.0625,0,0,0,0.375,0,0,0.0625,0,0.0625,0,0,0,0,0,0.0625,0,0,0.375,0.1875,0.0625,0.0625,0,0,0,0.0625,0.125,0,0.0625,0.0625,0,0.1875,0,0,0,0,0,0,0,0,0,0.125,0,0,0,0,0,0.6875,0.125,0.0625,0.4375,0,0.0625,0.625,0.0625,0.25,0,0,0,0,0,0,0,0.0625,0.1875,0,0,0,0,0.25,0.125,0.125,0.125,0.25,0.0625,0.125,0.1875,0,0.0625,0.1875,0,0,0.0625,0.125,0.0625,0,0,0,0,0.3125,0,0,0,0,0,0,0,0,0,0.0625,0.125,0,0,0.0625,0.0625,0,0.0625,0.3125,0.0625,0.3125,0.6875,0.125,0.5625,0.3125,0.0625,0.3125,0,0.0625,0,0.125,0.0625,0.25,0,0,0.0625,0,0,0,0.1875,0,0,0.0625,0.0625,0.0625,0.4375,0.375,0.4375,0,0,0,0.0625,0.0625,0.0625,0,0,0,0.3125,0.125,0.3125,0.1875,0.0625,0.125,0.125,0,0.125,0.5625,0.3125,0.375,0.4375,0.125,0.375,0.4375,0.3125,0.5,0.4375,0.25,0.375,0.3125,0,0.1875,0,0,0,0,0,0.125,0,0,0.0625,0,0,0,0,0.125,0,0,0.25,0.1875,0.4375,0.1875,0.5,0.4375,0,0.625,0.5625,0.0625,0.375,0.6875,0.1875,0.375,0,0,0,0,0,0,0,0,0,0,0,0.5625,0.0625,0.1875,0.4375,0,0.1875,0.125,0.375,0.375,0.6875,0,0.0625,0.25,0.125,0.125,0.125,0.6875,0.4375,0.75,0.5625,0,0.5,0.375,0.0625,0.125,0,0,0,0,0,0,0.25,0.3125,0.125,0,0,0,0,0,0,0,0,0,0.0625,0.1875,0.5625,0,0,0,0,0,0,0.1875,0.0625,0.3125,0.0625,0,0.125,0,0,0,0.3125,0.375,0.8125,0.4375,0,0.5,0,0,0,0.125,0.0625,0,0.0625,0.1875,0,0.3125,0.25,0.25,0.125,0.125,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0.0625,0,0.0625,0.125,0,0,0,0,0,0,0,0,0,0,0,0,0.125,0,0,0,0.25,0,0,0,0,0,0,0.125,0,0,0.0625,0.1875,0,0.125,0.1875,0.25,0,0,0,0,0,0,0,0,0,0.3125,0.4375,0.375,0.25,0.125,0.5625,0.375,0.125,0.4375,0.3125,0.1875,0,0.1875,0.125,0,0.5,0.0625,0.125,0.8125,0.5625,0.8125,1.25,0.1875,0.6875,0.0625,0,0,0.125,0,0,0.125,0,0,0.125,0,0,0,0.1875,0.375,0,0,0.25,0,0.1875,0.25,0.125,0,0,0.0625,0.125,0.0625,0.1875,0,0,0,0,0,0,0,0,0,0.125,0.0625,0,0,0,0,0,0,0.75,0.125,0.5,0,0.0625,0.0625,0,0,0,0,0,0,0.375,0,0.25,0.1875,0,0,0.75,0.375,0.5,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0.0625,0.0625,0.125,0,0,0,0,0,0,0,0,0,0.0625,0,0,0,0.0625,0,0.1875,0.1875,0.0625,0,0,0,0,0.0625,0.0625,0.125,0.25,0.4375,0.1875,0.0625,0,0.125,0,0,0,0,0,0.1875,0.1875,0.5625,0,0,0,0.3125,0.125,0,0,0.125,0,0.0625,0,0,0.125,0.125,0,0,0,0,0,0,0,0.1875,0.125,0.25,0.375,0.125,0.6875,0.375,0,0.125,0.3125,0.125,0,0.3125,0,0.1875,0.125,0.0625,0,0,0,0,0,0,0,0,0,0,0,0,0,0.125,0.0625,0,0,0,0,0.0625,0.1875,0.1875,0.125,0.1875,0.125,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0.1875,0.1875,0.1875,0,0,0.125,0.4375,0.1875,0.5,0,0,0,0,0.0625,0.125,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0.5,0.25,0.375,0.5,0.375,0.75,0.25,0.0625,0.75,0,0,0,0.1875,0,0,0.4375,0,0,0.3125,0,0,0,0,0.25,0,0,0,0.4375,0,0,0.375,0.125,0.0625,0,0,0,0,0,0,0,0,0,0.0625,0,0,0.1875,0,0,0,0,0,0,0,0.125,0.375,0,0,0,0.375,0,0.9375,1.4375,0.1875,0,0.3125,0,0,0,0,0,0.4375,0.875,0,0.5,0.5,0.4375,0.25,0.25,0,0.625,0,0.1875,0.1875,0,0,0,0,0,0,0,0.4375,0.0625,0.375,0.0625,0,0,0.5625,0,0.3125,0.25,0,0.125,0.125,0.375,0.5,0,0,0.3125,0.0625,0,0.5,0,0,0,0.5625,0.125,0.125,0.125,0.0625,0,0.125,0,0.6875,0,0,0,0.5625,0,0.1875,0,0,0,0,0,0,0,0,0.125,0,0,0,0,0,0,0.1875,1.125,0.25,0,0,0.0625,0,0,0,0,0,0.1875,0,0.3125,0,0.3125,1.375,0,0,0,0,0.3125,0,0,0.375,0,0,0,0,0,0.125,0.0625,0,0,0.1875,0,0,0,0,0,0,0,0.1875,0.25,0,0,0,0,0,0,0,0,0.3125,0,0.25,0.1875,0.1875,0,0,0,0,0,0,0,0.0625,0,0,0.0625,0.25,0.125,0.3125,0.625,0,0,0.375,0,0,0,0,0,0.125,0.25,0,0.1875,0.3125,0.1875,0.5,0.4375,0,0.75,0.5625,0,0,0.75,0.125,0.0625,0,0,0,0,0.125,0,0,0.875,0,0,0,0,0,0.0625,0,0.25,0.25,0,0,0,0,0.125,0,0.125,0.625,0,0.3125,1.0,0,0,0.1875,0,0,0,0,0.1875,0,0.125,0.75,0,0,0,0.375,0.0625,0.5,0.375,0,0.1875,0,0,0.0625,0,0,0,0,0,0.375,0,0,0,0,0,0,0,0.375,0.125,0,0,0,0,0,0,0.5625,0,0,0.375,0,0.0625,0,0,0,0,0.5,0,0,0,0,0,0,0,0.0625,0,0,0.1875,0,0.0625,0.3125,0,0,0,0,0,0,0.6875,0,0,0,0,0.3125,0.9375,1.5,0,0,0.1875,0.6875,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0.125,0,0.1875,0.0625,0,0,0,0,0,0.6875,0.3125,0,0,0,0,0.5,0.875,0.4375,0.3125,0.5,0,0,0.1875,0.6875,0.125,0.6875,0,0.25,0.5625,0.6875,0.1875,0.625,0.125,0,0.1875,0,0.125,0,0,0,0,0,0,0,0,0,0,0,1.125,0,0,0.75,0,0,0,0,0,0.0625,0,0,0,0,0,0,0,0,0.3125,0,0,0.0625,0,0,0,0,0,0.25,0,0,0,0,0,0,0,0.25,0.1875,0,0.375,0.8125,0.4375,0,0.25,0.0625,0,0,0,0,0,0,0.1875,0,0.25,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0.125,0.125,0,0.5625,0.0625,0,0,0,0,0,0.375,0.0625,0.5,0,0.1875,0,0,0,0,0.4375,0,0,0,0,0,0,0,0,0,0,0.875,0,0,0,0.375,0,0,0.1875,0.0625,0.0625,0.0625,0.125,0.25,0.75,0.25,0,0,0,0,0,0,0,0.4375,0.6875,0.625,0.6875,0.75,0,0,0,0,0,0,0.1875,0,0,0.375,0.75,0.1875,0,0.1875,0,0,0,0,0,0,0,0,0,0.125,0,0,0.125,0,0,0.0625,0.0625,0.9375,0,0,0.8125,0,0,0.4375,0,0.0625,0,0,0.8125,0,0,0.3125,0.25,0,0,0,0,0,0,0,0.25,0.25,0,0,0,0,0.5625,0,0.5,0.75,0,0.5625,0,0,0,0,0.0625,0,0,0,0,0.6875,0,0,0.1875,0,0,0,0.375,0,0.1875,0.4375,0.25,0,0,0,0,0.25,0,0.25,1.0625,0.1875,0.75,1.4375,0.5,0,0,0,0,0.1875,0.0625,0,0,0,0.1875,0.125,0.125,0,0,0,0,0,0.0625,0,0,0,0.125,0,0,0,0,0.125,0,0,0.0625,0,0,0,0,0,0,0.375,0,0,0.3125,1.3125,0.375,0,1.0,0,0,0.6875,0,0,0,0,0.0625,0,0,0.1875,0,0.125,0,0,0,0,0,0,0.0625,0.3125,0,0.125,0,0,0.5,0.8125,0.9375,0.8125,0.1875,0.8125,0.5,0.5,0.8125,0,0,0,0.8125,0,0.4375,0,0,0,0,0,0.125,0,0.5625,0.6875,0,0.3125,0,0,0,0.125,0,0.0625,0.3125,0.25,0.4375,0.5,0,0,0,0.1875,0,0.25,0,0,0,0.1875,0.1875,0,0,0.4375,0,0.375,0,0,0,0,0,0,0,0,0,0,0,0.75,0,0.4375,0.3125,0,0.125,0,0,0,0,0,0,0,0,0,0,0,0,0.125,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1.0,0.3125,0.75,0.9375,0,1.1875,1.1875,1.125,0.9375,0,0,0,0,1.4375,1.0625,0,0.0625,0.5,0.1875,0.125,0,0.0625,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0.5,0.625,0.25,1.0,0.5625,0,0.0625,0.25,0,0,0,0,0,0,0,0,0.5625,0.3125,0,0,0.1875,0,0,0,0,0,0,0,0,0,0.375,0,0.0625,0.25,0.4375,0.8125,0.9375,0.75,0.5625,0.125,0.375,0,0,0,0,0.8125,0,0,1.0625,0,0,0.9375,0,0,0,0.0625,0,0,0.1875,0.25,0,0,0.25,0,0,0,0,0,0,0.0625,0,0.4375,0,0.5,0.5625,0,0.8125,0.3125,0.125,0.25,0,0,0,0,0.9375,0,0,0,0,0.6875,0,0.6875,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0.25,0,0.375,0.75,0,0.4375,0,0.75,0,0.4375,0.875,0.5625,0,0,0.0625,0,0.0625,0.75,0,0,0,0.0625,0.1875,0,0,0,0,0.75,1.125,0.6875,0,0,0,0.125,0.3125,0,0.0625,0.0625,0,0.0625,0,0.125,0,0,0,0.4375,0,0.3125,0,0,0,0.4375,0.3125,1.0625,0,0,0.8125,0.5,0.0625,0.75,0.25,0.5,0.3125,0,0,0,0.125,0,0.25,0.1875,0,0,0.5625,0,0,0,0.8125,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0.125,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0.1875,0,0,0.4375,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0.25,0,0,0.125,0,0,0,0,0,0,0,0,0.5,0.25,0.4375,0,0.5625,0.625,0.375,1.3125,0.125,0.5625,0.6875,0.25,0,0,0,0.375,0.0625,0.125,0.375,0.1875,0.5625,0,0,0,0.5,0,0.8125,0.5,0.0625,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0.4375,0.3125,0.0625,0.625};

bias_s = '{0.03125,0.0078125,-0.1015625,0,0.21875,-0.015625,0.09375,0.3359375,0.15625,0,0.109375,0.1328125,0.0234375,-0.078125,-0.046875,0.0859375,0.03125,-0.0390625,0.078125,0.1328125,0.03125,0.03125,0.203125,-0.0625,0.09375,0,-0.0234375,0.0703125,-0.0703125,0.0078125,0.21875,0.0};

bias_1x1 = '{-0.015625,-0.015625,-0.046875,-0.015625,0,-0.0703125,0.0234375,-0.015625,-0.046875,0.015625,-0.03125,-0.0234375,-0.0390625,-0.015625,-0.078125,0.015625,-0.015625,-0.015625,0.03125,-0.0078125,0.0078125,-0.015625,-0.0390625,0.0078125,0.03125,-0.015625,-0.0234375,0.0234375,-0.015625,-0.0390625,0,-0.0078125,-0.03125,-0.03125,-0.0390625,-0.0234375,-0.0390625,-0.0078125,-0.015625,-0.0078125,-0.0234375,-0.0078125,-0.0078125,-0.046875,0.0078125,-0.03125,-0.015625,0,-0.015625,-0.0234375,-0.03125,-0.0390625,0,-0.03125,0,-0.0234375,-0.0234375,-0.0078125,0,-0.015625,-0.0625,0,-0.015625,-0.0390625,-0.0234375,-0.0078125,-0.0234375,-0.015625,0,-0.0078125,-0.03125,0.0234375,-0.015625,-0.09375,0.0078125,0.015625,-0.015625,-0.03125,-0.015625,-0.0546875,-0.0234375,-0.0390625,0.015625,-0.015625,0,-0.0078125,-0.0234375,0.0078125,-0.0078125,0,-0.03125,-0.1015625,-0.015625,-0.0234375,-0.0234375,0,-0.03125,-0.046875,-0.0078125,-0.03125,-0.015625,0,-0.015625,-0.046875,-0.046875,-0.0546875,-0.0546875,-0.0546875,-0.015625,-0.0234375,-0.0234375,-0.0078125,-0.03125,-0.015625,-0.015625,0.0078125,-0.03125,-0.0078125,-0.0859375,-0.015625,-0.0390625,-0.0234375,-0.0078125,-0.0234375,-0.0234375,0.015625,-0.046875,-0.0390625};

bias_3x3 = '{-0.015625,-0.046875,-0.0078125,0.0390625,0,-0.09375,-0.015625,-0.0546875,-0.015625,-0.09375,-0.0859375,-0.0234375,-0.015625,-0.0078125,-0.0390625,-0.03125,0.0234375,-0.0546875,-0.046875,-0.0234375,0.046875,-0.046875,-0.0390625,-0.0390625,-0.078125,0.0234375,-0.0703125,-0.046875,-0.1171875,-0.0546875,-0.0078125,0.0078125,-0.0390625,-0.0546875,-0.015625,-0.0078125,0,-0.0546875,-0.0546875,-0.046875,0,-0.0078125,-0.0234375,-0.0546875,-0.03125,-0.03125,0.0390625,-0.015625,-0.03125,-0.0234375,0.0078125,-0.0234375,-0.078125,-0.0625,-0.015625,-0.0234375,-0.0546875,-0.0703125,-0.0234375,-0.0546875,0.0078125,-0.0234375,-0.0234375,0,-0.0546875,0.015625,0.0234375,0.0078125,-0.0078125,0,0.046875,-0.046875,-0.0234375,-0.09375,-0.0703125,0.03125,0,-0.046875,-0.125,0.0078125,-0.1171875,0,0.0234375,-0.0234375,0.0078125,-0.03125,-0.0546875,0.0234375,-0.0703125,-0.0703125,-0.046875,-0.0625,0.0078125,-0.0390625,-0.0546875,-0.015625,0.0078125,0.03125,0,-0.0078125,-0.03125,-0.0390625,-0.0625,0.0390625,-0.015625,-0.0078125,-0.015625,-0.03125,0,0.0390625,0.078125,-0.1171875,-0.0625,-0.0625,-0.0546875,-0.0625,0,-0.046875,-0.046875,-0.03125,0.0234375,-0.015625,0.015625,0.0078125,0.015625,0.0234375,-0.015625,0.015625};

weight_s = '{-0.03125,0.0078125,0.03125,-0.015625,0,-0.0078125,0.0703125,-0.0234375,-0.03125,-0.0859375,0.0546875,-0.109375,-0.03125,0.0234375,0.03125,0.015625,0.0078125,-0.0390625,0,0,-0.0625,-0.0859375,0.046875,0,0.0390625,-0.0390625,-0.015625,0.03125,-0.0078125,-0.015625,-0.0390625,0.03125,0,0.0234375,0.03125,-0.015625,0.0078125,0,-0.0703125,0.0078125,-0.0234375,-0.03125,0.0078125,0.0859375,-0.0234375,-0.0078125,-0.078125,-0.109375,0.0234375,0.015625,0.046875,-0.046875,0.03125,0.0859375,-0.0078125,-0.0078125,0.0234375,0.015625,-0.0234375,0.0625,-0.1015625,-0.046875,0,-0.0390625,-0.0390625,-0.0390625,0.1171875,0.015625,-0.046875,0.0859375,-0.0390625,0.0078125,-0.015625,-0.078125,-0.0234375,-0.015625,-0.0546875,0.0078125,0,-0.0078125,-0.0234375,-0.0078125,0.1328125,0.0078125,-0.0234375,-0.0234375,-0.0078125,-0.0234375,-0.015625,0,-0.03125,-0.0234375,-0.0078125,0,0.0078125,0.015625,-0.078125,-0.0078125,-0.0625,-0.0703125,0.0546875,0.0390625,0.0546875,-0.0390625,-0.0078125,0.0078125,0.0703125,-0.046875,-0.0078125,0.046875,0.046875,-0.0390625,0.0078125,0.015625,-0.0390625,0.015625,0.0390625,0.0703125,-0.046875,0.015625,-0.0390625,-0.03125,0,-0.03125,-0.0703125,-0.0234375,-0.046875,-0.015625,-0.0703125,-0.1015625,-0.046875,-0.1171875,0.0859375,0.171875,-0.03125,-0.0625,0,0.1171875,0.125,-0.015625,-0.2265625,-0.015625,-0.09375,-0.1015625,0.109375,-0.0390625,-0.15625,0.03125,-0.0234375,0.015625,0.109375,-0.046875,-0.1796875,-0.0703125,0.0703125,-0.03125,0.0390625,0.0703125,-0.0390625,-0.1484375,-0.109375,-0.2109375,0.0234375,0.078125,-0.0234375,0.296875,0.0703125,-0.0390625,0.0625,-0.0703125,0.0625,0.03125,0.0625,-0.09375,0.140625,-0.1328125,0.0859375,0.140625,0.078125,0.03125,0.015625,-0.0625,0,0.078125,0.0703125,-0.109375,0.0859375,-0.078125,0.1171875,-0.0703125,-0.0625,-0.015625,-0.0546875,-0.0390625,-0.0703125,0.03125,-0.046875,-0.0234375,0.0234375,0.2421875,-0.0078125,-0.140625,-0.1640625,0.0390625,0.0078125,0.046875,-0.015625,0,-0.03125,0.046875,-0.09375,-0.0234375,0.0234375,0.0390625,0.0234375,-0.0078125,-0.046875,0.0234375,-0.015625,0.1328125,-0.0390625,-0.0234375,0.1171875,-0.0390625,0.109375,0.03125,0.203125,0.140625,-0.0625,-0.1328125,-0.046875,0,-0.0625,-0.0234375,0.140625,0.0703125,-0.078125,0,0.109375,0,-0.0078125,-0.0546875,0.1171875,0.03125,-0.1015625,0.1015625,-0.0390625,-0.109375,-0.0625,0.1328125,0.0859375,0.1640625,0.015625,-0.0234375,-0.078125,0.046875,0.0234375,0.0234375,0.0078125,-0.015625,-0.015625,-0.0078125,-0.0234375,0.03125,0.0234375,0.0625,-0.0078125,-0.015625,0.0078125,-0.015625,-0.015625,0.0078125,-0.0078125,-0.0078125,0,0.015625,0,0.015625,-0.0078125,0.0078125,0,0.0078125,-0.0078125,-0.0078125,0.0078125,-0.015625,0.0078125,-0.015625,0,0,0.0234375,0.03125,-0.0234375,-0.0234375,0.0234375,-0.0390625,0.0234375,0,0.0078125,-0.015625,0.015625,0.0078125,0,0.0234375,0.015625,0.015625,0.015625,0.015625,0.0078125,0.015625,0.015625,0,0.03125,0.0234375,0.015625,-0.0234375,0.03125,0.015625,0.0078125,0.015625,-0.0078125,0.0078125,0.015625,0.0078125,0.015625,0.0234375,-0.015625,0.0078125,-0.015625,0.015625,-0.015625,-0.0078125,-0.015625,0.0078125,0,0.015625,0.015625,0.015625,-0.015625,0,0.03125,0.015625,-0.0078125,-0.0234375,-0.0234375,-0.0234375,0.015625,0.0234375,-0.0078125,0.0078125,0.0078125,-0.015625,0.0390625,0,0.0078125,0.015625,-0.0390625,0.0078125,-0.015625,0.0078125,0,-0.0078125,-0.015625,-0.015625,0,0.015625,-0.0078125,-0.0078125,-0.0078125,0.015625,0,0.015625,0,0,0,-0.0078125,0.0078125,0,0.015625,0,0.015625,0.015625,0,-0.0078125,0,-0.0078125,-0.0078125,0,0.015625,0,0.015625,-0.0078125,-0.0234375,-0.0078125,-0.0078125,-0.0234375,-0.0078125,0,0,0.0078125,-0.0234375,0.015625,0.015625,0.0078125,0,0.0078125,-0.0234375,-0.0234375,-0.0234375,-0.03125,0.015625,-0.0078125,-0.015625,0.03125,-0.0234375,-0.03125,-0.0078125,0,0.0078125,0,0,0.0078125,-0.03125,0.03125,0.0234375,0.015625,0.015625,0.0234375,0,0.0234375,0.015625,-0.015625,0.0078125,-0.0078125,0,-0.015625,0.0078125,-0.0078125,0.015625,0.03125,0,-0.015625,-0.015625,-0.015625,-0.0078125,-0.015625,-0.0078125,0.015625,-0.03125,0.0078125,-0.0234375,0.0234375,0.0078125,0.015625,-0.0078125,-0.015625,0.015625,0.0078125,-0.0078125,-0.015625,-0.0234375,-0.0078125,-0.0234375,0.0234375,0.0078125,-0.0078125,0.015625,0.0234375,0.0234375,0.0078125,0.03125,-0.0078125,-0.015625,-0.0078125,-0.0625,0.015625,0,0.015625,-0.0078125,0.0234375,-0.0078125,0,0.0078125,0.015625,-0.0234375,-0.0234375,-0.0078125,0.046875,-0.0078125,-0.015625,-0.03125,-0.015625,-0.015625,0,0.0078125,0,-0.0078125,-0.0078125,0.03125,0,0.0078125,0,0,0,-0.0234375,-0.0078125,-0.0390625,-0.0234375,-0.015625,-0.0078125,0.015625,-0.0078125,0.0859375,0.078125,0.0078125,0.046875,-0.0234375,-0.0078125,0,0.1171875,-0.0078125,-0.1328125,-0.0625,-0.0078125,0,-0.046875,0.0078125,0,0,0.0703125,-0.0078125,0.046875,0.015625,0.0390625,0.109375,-0.03125,-0.0390625,0.1015625,0.0234375,-0.0390625,0.0078125,0.015625,0.015625,-0.0078125,-0.015625,0.1171875,0.0546875,0,-0.0078125,0.1328125,-0.0546875,0.0390625,-0.03125,0.03125,-0.03125,0.078125,0.046875,0.0234375,0.1640625,0.03125,0.015625,0.0546875,-0.1015625,0.046875,-0.0078125,0.0390625,0.0390625,0.0078125,0.0546875,-0.0546875,0.0390625,0.0078125,0,0.0078125,-0.0234375,-0.015625,0.015625,0.0078125,-0.0546875,0.0234375,-0.046875,-0.0078125,-0.0234375,0.046875,0.0703125,-0.03125,0.03125,-0.03125,-0.0078125,0.046875,0.0625,-0.0390625,0.0546875,0,0.15625,0.0703125,0.09375,-0.03125,-0.0078125,0.046875,0.03125,0.140625,-0.0078125,-0.015625,0.0234375,0.015625,0.015625,0.125,0,0.03125,0.0625,-0.046875,0.0390625,-0.0078125,0.0703125,0.0234375,-0.0078125,-0.0546875,0.0234375,-0.0234375,-0.0078125,-0.078125,0.0078125,-0.015625,-0.015625,0.0390625,0.0625,0.0234375,0.0234375,0.0625,0.0078125,-0.0078125,0,0.09375,0,-0.03125,0.0546875,-0.046875,-0.0625,0.0703125,0.078125,0.0859375,-0.0390625,-0.0859375,0.1171875,0.0703125,-0.0234375,0.0390625,-0.046875,-0.0390625,-0.046875,-0.0546875,-0.125,-0.0390625,-0.0703125,-0.046875,0.0078125,0.0078125,-0.03125,0.015625,-0.0859375,0.0390625,0.125,0.078125,0.09375,0.0234375,0.0390625,-0.0078125,0.140625,-0.0390625,-0.09375,-0.09375,-0.109375,-0.1796875,0.046875,0.0078125,0.015625,-0.015625,0.109375,0.078125,-0.0703125,0.0546875,-0.0703125,-0.0234375,0.0390625,-0.0546875,0.1640625,-0.03125,-0.0625,0.0390625,-0.109375,-0.046875,0.0390625,0.046875,0.015625,-0.0625,-0.0390625,0.0390625,-0.0703125,0.015625,0,0.0390625,0,0.09375,0.0234375,-0.0546875,-0.0546875,-0.1015625,0.015625,0.015625,0.0625,0.078125,-0.0234375,0.0390625,-0.03125,-0.0703125,-0.046875,-0.0390625,0.0078125,-0.1640625,-0.0234375,-0.0390625,-0.1015625,0.0078125,-0.1015625,-0.0859375,-0.0625,0.03125,0.140625,0.1015625,0.015625,0.203125,0.09375,-0.078125,0.1171875,0.046875,-0.171875,0.0703125,0.0078125,0.2421875,-0.015625,-0.109375,-0.046875,-0.0625,0.0546875,0.0546875,-0.0703125,-0.0078125,0.1015625,-0.046875,0,0.046875,0.0625,0.09375,-0.09375,-0.0078125,0.0546875,0.0234375,-0.0234375,-0.140625,0.015625,0.015625,-0.03125,-0.0234375,-0.015625,0.0859375,0.109375,-0.0234375,0.0390625,0.03125,-0.0546875,0,0.0078125,0.0078125,-0.0390625,-0.09375,-0.0234375,-0.03125,0.015625,-0.0390625,-0.0078125,0.0859375,0.015625,-0.015625,0.0078125,-0.0234375,0.015625,0.0078125,-0.0625,-0.03125,-0.03125,0,0.0625,0.0546875,0.0078125,0.046875,0.0234375,-0.0390625,0.0625,0.046875,-0.0234375,0.0234375,-0.0234375,-0.0546875,0,0.0078125,-0.0390625,0.1640625,-0.03125,0.015625,0.0859375,0.0546875,0.015625,0.0703125,0.0546875,0.03125,0.0234375,-0.0078125,-0.0390625,-0.0078125,0.1015625,-0.09375,-0.015625,-0.0390625,0.03125,-0.0078125,0.0859375,0.0625,-0.0078125,0.046875,-0.015625,-0.0390625,-0.078125,-0.0546875,-0.0546875,0,-0.0390625,-0.015625,0,0.109375,-0.0390625,0.0625,0.046875,-0.03125,0.0390625,0.03125,0.03125,-0.0234375,0,0,0.0625,0.0078125,0.0234375,0.0703125,-0.0078125,-0.0078125,0.0234375,-0.015625,-0.0390625,-0.0234375,-0.0078125,0,0.03125,0.0078125,-0.03125,-0.015625,0.0078125,-0.03125,0.03125,-0.0390625,0.0390625,-0.0234375,-0.03125,-0.046875,-0.0078125,-0.015625,-0.0078125,-0.015625,-0.03125,0,0.015625,0.0234375,0.0078125,-0.0234375,-0.0078125,0.03125,-0.0625,-0.0078125,-0.0234375,0.0234375,0.0078125,-0.0390625,0.0078125,0.015625,-0.0625,0.0234375,-0.0234375,0.2890625,-0.0625,-0.0234375,-0.0703125,0.0703125,-0.0234375,-0.03125,-0.15625,-0.0234375,0.0078125,-0.0078125,-0.0625,-0.015625,0.125,-0.140625,-0.1015625,0.0390625,0,0.109375,-0.0390625,-0.046875,-0.03125,0.0390625,0.078125,0.09375,-0.015625,0.0234375,0.0078125,-0.03125,0.140625,0.0859375,-0.03125,-0.1171875,-0.125,-0.0625,0.0390625,0.015625,0.1640625,0.0390625,-0.03125,-0.09375,0.015625,-0.03125,0.1171875,0,-0.0625,0.0078125,-0.0078125,-0.078125,-0.0390625,0.0078125,-0.0390625,-0.0859375,-0.078125,0.0859375,-0.015625,0.0625,-0.0234375,-0.0390625,-0.03125,0.0625,-0.1328125,0.0234375,-0.015625,-0.0234375,0.0078125,-0.015625,-0.09375,0.046875,-0.1171875,-0.0546875,-0.0546875,0.125,0.2109375,0.1796875,-0.078125,-0.0078125,0.046875,-0.0859375,-0.0859375,-0.046875,0,-0.0625,-0.015625,0.1015625,0.03125,-0.09375,-0.09375,-0.0234375,-0.1171875,-0.0390625,0.0625,-0.0703125,0.015625,-0.109375,-0.109375,-0.0234375,0,0.0234375,0.1015625,0.078125,0.109375,0,0.0703125,-0.0703125,0.171875,-0.03125,0.125,0.0078125,-0.046875,0.1015625,-0.0078125,-0.0703125,0.0234375,-0.0078125,-0.046875,0.0625,0.0546875,0.03125,-0.0234375,0.0078125,0.046875,0.0234375,-0.0078125,0.0859375,0.15625,-0.09375,-0.03125,0.046875,-0.03125,0,-0.0078125,0,-0.0078125,0.0859375,0.0390625,-0.0234375,-0.0546875,-0.0859375,-0.0078125,0.0234375,-0.0390625,-0.015625,-0.0078125,0.1484375,-0.0390625,-0.0390625,0.0234375,0,-0.0078125,0.0390625,-0.1171875,-0.0625,0.0546875,-0.03125,-0.0546875,-0.0234375,-0.0625,-0.0078125,0.0078125,0,-0.0390625,0.0390625,0.015625,0,-0.03125,-0.0703125,0.015625,0.0078125,-0.0078125,0.0078125,-0.0234375,-0.03125,0,-0.0234375,-0.0078125,-0.0078125,0,0.015625,-0.046875,0.0546875,-0.015625,0.0234375,0.046875,0,-0.1171875,-0.0390625,-0.03125,-0.0859375,-0.0234375,0.0234375,-0.03125,0.0234375,0.0546875,0.015625,0,-0.0859375,-0.0546875,0.0546875,0.0390625,0.03125,-0.0078125,-0.046875,-0.078125,0.1171875,0.0078125,0.0078125,-0.015625,0.015625,-0.015625,-0.015625,-0.0625,0.0234375,0,-0.0078125,0.0078125,0.0390625,0.0078125,-0.0390625,0.0078125,-0.015625,-0.0234375,0.0234375,0.125,0.015625,0.03125,0.0859375,0.0234375,-0.015625,-0.0234375,0.0078125,0.0234375,-0.0390625,0.0078125,-0.0625,-0.0078125,-0.1015625,-0.0234375,0.015625,-0.0078125,0.0625,-0.046875,-0.015625,-0.015625,-0.03125,0.03125,-0.015625,-0.0546875,-0.0234375,0.015625,-0.0390625,0.0625,-0.03125,0.015625,-0.0390625,0.0234375,-0.1328125,0.0390625,-0.0234375,-0.0625,0.015625,-0.1875,0.0390625,0.1171875,0.203125,-0.03125,0.046875,-0.1953125,0.0078125,-0.140625,0.0859375,-0.0703125,0.0546875,0.2265625,0.171875,0.0703125,-0.0234375,-0.234375,0.0390625,-0.015625,0.0390625,-0.0078125,0.0078125,0.0078125,0.0703125,0.015625,0.0078125,-0.15625,0.03125,0.0078125,0.046875,-0.015625,0.0546875,-0.1640625,0.1640625,-0.03125,-0.125,0.3046875,-0.015625,-0.0625,0.0390625,-0.0625,-0.1640625,-0.09375,0.078125,0,0.09375,0.0859375,-0.1015625,-0.0859375,-0.046875,0.0546875,-0.015625,-0.03125,-0.09375,-0.1796875,-0.078125,0,0.0078125,-0.09375,0.109375,0.0546875,-0.15625,0.140625,-0.0625,-0.03125,0.0234375,-0.078125,0.015625,-0.046875,0.1328125,0.09375,0,-0.1484375,0.078125,-0.09375,-0.09375,-0.0625,-0.1015625,0.0703125,-0.0625,-0.1328125,-0.109375,-0.015625,0.09375,-0.078125,-0.0078125,0.078125,-0.0859375,-0.1171875,0.0546875,0.1171875,-0.03125,0.0234375,0.0625,0.0390625,0.1171875,-0.046875,0.0078125,0.0078125,-0.1171875,-0.0234375,0.0234375,0.0546875,-0.0859375,0.03125,0.0859375,0.09375,-0.1171875,0.0703125,0.2109375,0.1875,0.015625,0,0,-0.0078125,-0.1328125,-0.140625,-0.140625,0.046875,0.109375,0.1015625,-0.0625,-0.0234375,-0.0078125,-0.015625,0.0078125,0,0.0078125,-0.0078125,0,-0.0078125,-0.0078125,0.015625,0.0078125,0,-0.0234375,-0.0234375,0.015625,-0.015625,-0.015625,-0.0078125,0,0,-0.015625,-0.015625,0.015625,0,-0.015625,0,0,0.0078125,-0.0078125,0.0078125,-0.0078125,-0.0078125,-0.015625,0,0.0078125,0,0,-0.0078125,-0.015625,0.015625,-0.015625,-0.0078125,-0.0078125,0,0.0078125,-0.0078125,0,0.0078125,-0.0078125,0,-0.015625,0,-0.0078125,-0.0078125,0,0,-0.0078125,0.0078125,0.0078125,-0.015625,-0.015625,0,0,-0.0078125,-0.0078125,-0.0078125,0.0078125,-0.015625,0.015625,0.0078125,-0.0078125,-0.015625,-0.015625,-0.0078125,0,-0.0078125,-0.015625,-0.0078125,0,0,0,-0.015625,-0.015625,-0.0234375,-0.0078125,0,0,-0.015625,-0.015625,0.0078125,-0.0078125,0.0078125,0,-0.0078125,-0.0078125,-0.0234375,-0.015625,0,-0.0078125,0.015625,0,-0.0078125,0,-0.0078125,-0.0078125,-0.0078125,0,-0.0078125,-0.0078125,0,0.0078125,0,-0.0078125,0,-0.0078125,0.0078125,0,0.0078125,-0.0078125,0,-0.015625,0,-0.015625,-0.0078125,0,-0.015625,-0.015625,-0.015625,0.0078125,0.0078125,-0.015625,-0.015625,0.0078125,-0.015625,-0.0234375,0.0078125,0,0.0078125,0,0,0.015625,-0.0078125,0,-0.0078125,-0.015625,0,-0.0078125,-0.0078125,-0.015625,-0.015625,0.0078125,0,-0.0078125,0.015625,-0.0078125,0,-0.0234375,0,-0.015625,0.015625,0.0078125,0.0078125,-0.0078125,0.0078125,0,0.0078125,0.0234375,0.0078125,0,-0.015625,-0.0234375,0.0234375,0,0.015625,0.0078125,0.015625,0.0078125,0,-0.0078125,0,-0.0078125,-0.0078125,-0.0234375,0,0.0078125,0.015625,0.0078125,0.0078125,0,-0.0078125,-0.0078125,0,0,0.0078125,-0.015625,0.0078125,0.0078125,0.0078125,-0.015625,-0.0078125,-0.015625,0.015625,-0.015625,-0.015625,0,-0.0078125,0.0078125,0.015625,-0.015625,0.0078125,0.0078125,-0.0078125,-0.015625,-0.015625,0.0234375,0.03125,0.015625,-0.015625,0.0234375,0.015625,-0.015625,-0.0078125,0,-0.0078125,-0.0234375,-0.015625,0.0546875,-0.0078125,-0.0078125,0.015625,0,0.015625,-0.0078125,-0.015625,0.015625,-0.0078125,0.0078125,0,0,-0.0078125,0,0.03125,0.0078125,0.015625,0.03125,0.0078125,0,0,-0.0078125,0,0.03125,-0.0078125,-0.015625,-0.0078125,0.0078125,0.078125,0.1171875,0.046875,0,-0.03125,0.0078125,-0.015625,0.078125,0.015625,0.046875,-0.09375,-0.09375,-0.046875,-0.0625,0.0703125,0,0,0.078125,-0.046875,-0.0390625,0.0078125,-0.0703125,-0.0546875,-0.015625,0.0078125,0.015625,0.046875,0.015625,0.0625,0.0078125,0.0078125,-0.03125,-0.0078125,-0.0078125,0.0078125,0.078125,0.109375,-0.0546875,0.03125,-0.0546875,0.140625,-0.0078125,0.015625,0.125,0.1328125,-0.0390625,0.015625,-0.015625,-0.0390625,0.0859375,-0.0234375,0.0234375,0.0546875,0.0625,0.046875,0.015625,0.0546875,-0.03125,0.0390625,-0.0703125,0.046875,0.046875,-0.0078125,0.015625,-0.0703125,0,-0.046875,0,0.15625,-0.0078125,-0.0078125,0.0078125,-0.015625,0.1015625,0.046875,-0.078125,-0.0703125,-0.0078125,0.0078125,-0.03125,0.0078125,0.03125,-0.015625,-0.0078125,-0.03125,-0.0546875,-0.0078125,0.0078125,0.015625,-0.046875,-0.015625,0.0078125,-0.046875,0.015625,0.09375,-0.03125,-0.0078125,-0.0390625,0.046875,0.015625,-0.046875,-0.0390625,-0.015625,0.125,0.0390625,0.0234375,0.0625,-0.0625,0,-0.046875,-0.03125,-0.0390625,0.03125,0.15625,0.0390625,0.0234375,0.015625,0.0390625,-0.0390625,0,-0.0234375,0.046875,0,-0.125,0.1328125,0.03125,-0.03125,-0.0390625,0.09375,0.0859375,0.1875,-0.046875,0.015625,-0.0234375,0.0703125,-0.1328125,-0.0234375,0.0234375,-0.15625,-0.171875,0.0078125,-0.0234375,-0.1015625,-0.078125,-0.0234375,-0.0703125,0,0.0546875,0.0703125,-0.03125,0.078125,-0.0390625,0.0078125,0.0390625,0,0.03125,0.03125,-0.09375,0.0859375,0.1875,-0.1015625,0.0390625,-0.1328125,-0.0390625,0.046875,-0.0625,0.2109375,-0.140625,0.09375,-0.0078125,-0.03125,-0.03125,-0.0546875,0.03125,-0.015625,-0.046875,-0.0625,-0.0625,-0.0390625,0.078125,-0.0078125,-0.171875,0.0625,0.171875,-0.1171875,-0.03125,-0.0546875,0.0078125,-0.0390625,-0.015625,-0.1171875,0,0.0546875,-0.015625,0.1328125,-0.0390625,-0.0703125,0.0859375,0.09375,0.0234375,-0.015625,0.109375,-0.0859375,0.0390625,-0.046875,0,-0.078125,0.140625,-0.0859375,-0.1015625,-0.0390625,0.015625,-0.140625,0.1015625,-0.015625,-0.09375,0.015625,-0.0703125,0.0390625,0.0078125,-0.0546875,-0.015625,-0.0546875,0.1875,0.0234375,0.1015625,-0.15625,0.0625,0.0234375,-0.1484375,-0.09375,-0.09375,0.15625,-0.140625,-0.109375,0.09375,0.0234375,-0.0859375,-0.1015625,-0.078125,-0.1953125,-0.0703125,0.0234375,0.0234375,-0.03125,-0.1171875,0.0390625,0.171875,-0.0703125,-0.0546875,-0.0703125,-0.078125,0.03125,-0.015625,-0.1015625,0.078125,0.0546875,0.015625,0.078125,-0.015625,-0.0234375,0.0078125,-0.0625,0.0546875,0.015625,-0.078125,-0.078125,0.0546875,-0.046875,0.0625,0,0.0546875,0.0078125,0.078125,0.0078125,-0.0234375,-0.0234375,-0.0078125,-0.0078125,0.109375,-0.0078125,-0.046875,-0.015625,0,-0.0234375,0.03125,0.1015625,0,0.015625,0.09375,0.015625,0.015625,-0.046875,-0.0546875,0.078125,0.03125,-0.015625,0.046875,-0.0390625,0,-0.015625,-0.09375,-0.015625,-0.0859375,-0.078125,-0.0234375,0.03125,-0.015625,-0.0546875,-0.0234375,-0.0078125,0,0.0703125,0.03125,-0.0078125,0.015625,0.0390625,0.015625,0,-0.015625,-0.0625,0.0234375,0.0234375,0.0078125,-0.0078125,0.015625,0.0078125,-0.0703125,0,-0.0234375,0.015625,-0.0390625,-0.1328125,-0.15625,0.046875,0.0859375,-0.1484375,-0.03125,0.0546875,0.0078125,-0.0546875,0.0078125,0,-0.0078125,-0.03125,-0.0234375,0.015625,0.0625,0.03125,-0.0078125,-0.046875,0.03125,0.03125,-0.0546875,-0.0546875,0.1015625,-0.0859375,-0.0546875,0.0234375,0.0546875,-0.078125,0.0390625,0.0546875,-0.1328125,0,0.046875,0.0078125,-0.0078125,0.0546875,-0.0859375,-0.0546875,-0.03125,-0.0625,-0.140625,-0.015625,-0.0078125,-0.0625,-0.0859375,0,-0.0390625,-0.0859375,-0.0703125,-0.0390625,-0.1015625,-0.046875,-0.1171875,-0.0703125,0.125,0.1640625,0.03125,-0.1015625,0.203125,0.1015625,0.0625,0.1484375,-0.0859375,-0.046875,0.1875,0.015625,0.015625,0.0078125,-0.1640625,-0.0234375,-0.0625,0.046875,0.1328125,-0.1015625,0.0703125,0.1953125,0.015625,-0.0078125,0.1640625,-0.0625,0.0859375,0.1328125,-0.171875,0.09375,0,0.0703125,0.0234375,-0.078125,0.0390625,0.1328125,-0.0078125,-0.109375,0.109375,0.046875,-0.1328125,0.0234375,-0.0390625,-0.09375,-0.078125,0.109375,0.1640625,-0.140625,0.109375,0.0859375,0.0546875,-0.1328125,-0.0546875,0.0625,0.03125,-0.015625,-0.0859375,-0.0859375,-0.0078125,-0.078125,0.03125,-0.0859375,0.046875,-0.078125,-0.0078125,0.0078125,0.078125,-0.0234375,0.140625,0.078125,-0.0703125,0,-0.1171875,-0.171875,0.2578125,0.0703125,-0.0703125,-0.0390625,-0.046875,-0.0546875,0.03125,-0.1328125,0.015625,-0.203125,0.1328125,-0.03125,-0.0078125,-0.1953125,-0.1328125,0.03125,0.2421875,0.078125,-0.0703125,-0.109375,-0.0078125,-0.0546875,-0.140625,0.0390625,-0.140625,-0.0703125,-0.0546875,0.0390625,0,0.0625,-0.1171875,0.03125,0.203125,0.1171875,0.1640625,-0.109375,0.0625,-0.0234375,0.125,-0.0625,0.0078125,-0.1015625,0.03125,0.125,-0.0625,-0.0234375,0.15625,0.078125,0,-0.0078125,0.0390625,-0.0546875,-0.0390625,0.0234375,0,0,0,-0.0390625,0.046875,-0.015625,-0.0390625,0.0390625,0.046875,0.0078125,0.140625,0.0234375,0.0078125,-0.0078125,0.0859375,0.09375,-0.0078125,-0.0625,0.0390625,0.0234375,-0.0234375,0.03125,-0.0390625,0.0078125,0.0625,0.1015625,0.0078125,-0.046875,0.0234375,0.0078125,-0.015625,-0.03125,0.0546875,-0.015625,-0.015625,0.015625,0.1171875,0.015625,-0.015625,-0.0078125,0.1171875,-0.046875,-0.109375,0.03125,0.0078125,0.015625,0.0546875,0.09375,-0.0546875,0.0546875,0.0703125,0.0390625,0.03125,0.0234375,0.0625,0.0390625,0.0546875,-0.03125,-0.0390625,0,0,-0.046875,-0.078125,0,-0.0078125,-0.0078125,0,-0.015625,-0.0078125,0.1171875,-0.015625,0.0078125,0.03125,-0.0390625,0.015625,0.03125,-0.015625,-0.0234375,0,0.015625,-0.015625,-0.015625,-0.109375,0.0078125,0.078125,0.0078125,0.0703125,-0.0546875,-0.0390625,-0.0078125,-0.015625,0.03125,0.1015625,0,-0.015625,-0.0390625,-0.015625,-0.1484375,-0.0234375,0.0390625,-0.0703125,-0.0078125,0.015625,0.03125,0.0078125,-0.0078125,0,-0.015625,0.0078125,-0.03125,-0.0625,0.0078125,0,0.1328125,-0.0078125,0.078125,0.015625,0.015625,-0.0234375,-0.0078125,-0.0703125,0,-0.015625,-0.0546875,-0.1171875,-0.078125,0.0625,0.234375,0.046875,-0.0234375,-0.09375,-0.1796875,0.0234375,0.0390625,0.09375,0.0546875,-0.078125,-0.1171875,0.0546875,-0.078125,-0.015625,-0.109375,-0.0078125,0.0234375,-0.078125,-0.03125,0.1484375,0.09375,-0.2109375,-0.0703125,0,-0.1015625,0.0078125,0.0703125,-0.0546875,0.140625,-0.0390625,0,0.1328125,0.1796875,-0.03125,0.046875,-0.09375,0.0078125,0.078125,-0.0546875,-0.1015625,0,-0.203125,0.1171875,0.125,0.0625,-0.1015625,-0.140625,0.0703125,0.0234375,0.1015625,0.109375,0.0234375,-0.1328125,-0.046875,0.1484375,0.03125,0.0546875,-0.015625,0.046875,0.0546875,0.046875,0.171875,-0.1171875,-0.0859375,-0.0234375,-0.0625,0.125,-0.140625,-0.1953125,-0.0078125,-0.0625,0.0234375,0.09375,-0.0078125,0.0234375,-0.109375,-0.09375,-0.1015625,-0.2890625,-0.0625,-0.03125,0.03125,-0.1484375,0.078125,-0.171875,-0.015625,0.1328125,0.09375,-0.15625,-0.046875,0.09375,0.03125,-0.09375,-0.015625,0.1328125,0.2265625,0.1640625,0.03125,0.078125,0.0390625,0.046875,0.0546875,-0.015625,-0.109375,0.140625,-0.2265625,-0.0625,-0.1796875,0.1953125,0.0546875,0.046875,-0.109375,-0.1640625,0.0234375,0.0390625,-0.140625,0.1796875,0.015625,-0.109375,0.0234375,-0.03125,-0.1328125,-0.0546875,-0.1171875,0.046875,-0.0703125,0.0078125,-0.03125,-0.0234375,-0.03125,0.046875,0.015625,0.015625,-0.0390625,-0.0234375,-0.0625,0.0390625,0.03125,0.0546875,-0.046875,-0.015625,-0.015625,0.0078125,-0.0625,0.0078125,0.0390625,0.0703125,0.09375,0.1796875,-0.0625,-0.0390625,-0.0078125,0.046875,0,0.0234375,0.0234375,-0.078125,0.046875,-0.015625,0,0,0.015625,0.015625,0.1171875,-0.03125,-0.1015625,-0.0546875,0.0546875,-0.109375,0.015625,-0.0390625,0.0390625,-0.0703125,-0.0390625,-0.0234375,0.0625,-0.03125,0.015625,-0.0078125,0.015625,0,-0.0078125,-0.0078125,-0.03125,-0.0234375,0.03125,-0.03125,0,0.0078125,0.03125,-0.03125,0.1015625,-0.0078125,-0.0234375,0.015625,0.0546875,-0.015625,-0.0546875,0.015625,0.0390625,0.0078125,-0.0234375,-0.0390625,-0.0234375,0.0078125,-0.0390625,-0.0078125,0.0234375,0.125,-0.03125,0.03125,0.015625,0,0.1015625,0.0078125,0.078125,-0.0625,-0.03125,0.0234375,0,0.0390625,0.109375,0,0.125,-0.015625,-0.1171875,0.078125,0.0078125,0,0.03125,0.0625,-0.0625,0.015625,0.015625,0,0.0234375,0.0078125,0.046875,0.0546875,-0.0859375,0.0390625,0.078125,-0.0390625,0.03125,0.0390625,0.015625,0.015625,-0.0078125,0.0078125,0.0390625,0.0234375,-0.03125,0.015625,-0.0234375,0.1171875,0.0703125,-0.015625,0.015625,0.1015625,0.015625,0.0078125,-0.0078125,-0.0703125,-0.0078125,-0.03125,-0.0078125,0.0234375,0.109375,0.078125,0.0234375,0.015625,-0.015625,-0.1171875,0.015625,-0.0703125,0.078125,0.125,-0.03125,-0.0546875,0.046875,0.0703125,0.0859375,-0.015625,0.0390625,-0.0546875,-0.0390625,0.1015625,0.015625,-0.015625,0.0703125,0.0546875,0,0.03125,-0.015625,-0.046875,0,0.015625,-0.0234375,0.0234375,-0.0234375,0.09375,0,-0.0859375,-0.046875,-0.0390625,-0.0703125,-0.0078125,0.109375,0.046875,-0.0546875,0.0390625,-0.03125,0.078125,-0.0078125,0.0078125,0,-0.0703125,-0.046875,-0.09375,0.0078125,-0.09375,-0.0234375,-0.015625,-0.078125,0.015625,0.03125,0.03125,0.1015625,-0.0390625,-0.0859375,-0.1328125,0.046875,0.03125,-0.015625,0.0625,0.078125,0.03125,-0.0390625,-0.0625,-0.0234375,-0.0390625,0.078125,0.03125,0.109375,0.09375,-0.0234375,-0.0390625,0.0390625,0.1328125,0.109375,-0.046875,-0.03125,-0.1171875,-0.0390625,-0.015625,-0.015625,-0.0546875,-0.015625,0.0078125,0.015625,-0.109375,-0.0390625,-0.03125,-0.0390625,-0.0234375,-0.0078125,-0.03125,-0.0703125,0.0234375,0.03125,-0.09375,0.03125,0.0859375,-0.078125,0.1484375,0.1015625,-0.09375,0.0390625,-0.0390625,-0.046875,0.03125,-0.0234375,-0.0078125,-0.03125,0.0234375,-0.015625,-0.0625,0,-0.0703125,0.0703125,0.015625,0.0859375,-0.0234375,-0.03125,-0.0390625,-0.015625,0.015625,-0.015625,-0.0078125,0.046875,-0.03125,-0.015625,-0.046875,0.015625,-0.09375,0.0234375,-0.0234375,0.03125,-0.046875,-0.0078125,0.0546875,-0.0234375,-0.0078125,-0.0234375,0.0078125,0.0625,0.0546875,0.03125,-0.0859375,-0.0703125,0.0859375,0.0234375,0.09375,-0.015625,0,0.09375,0,-0.0625,-0.015625,0.03125,-0.0234375,0.0703125,0.15625,-0.03125,0.1484375,0.0078125,0.0078125,0.046875,-0.0078125,0,-0.0546875,-0.0859375,0.1640625,-0.046875,0.0234375,0.046875,-0.1875,-0.0234375,0.0859375,-0.015625,-0.0234375,0.0078125,0.0234375,-0.0546875,-0.0234375,0.0625,-0.0078125,-0.0390625,0.0078125,0.015625,-0.0078125,0,0.03125,0.0078125,-0.0703125,0,-0.0390625,0.015625,0,-0.0703125,-0.046875,-0.03125,0.0546875,-0.015625,-0.0078125,0.0078125,0.1171875,0.0078125,0.015625,-0.09375,0.015625,-0.03125,-0.203125,-0.046875,0.09375,-0.0625,0.0703125,0.1015625,-0.0078125,0.1015625,-0.0078125,0.0703125,0.015625,0,0.1171875,0.015625,0.015625,-0.078125,0.15625,-0.0234375,-0.0234375,-0.015625,0.0703125,0.0234375,0,0.015625,-0.1015625,0.0234375,0.0234375,-0.1171875,-0.015625,0.03125,0.0234375,-0.109375,-0.0625,-0.0546875,-0.078125,-0.0078125,0.1796875,-0.0546875,0.09375,0,-0.0234375,0.078125,-0.1171875,0,0.046875,0.03125,0.046875,-0.03125,0.140625,0.0703125,-0.0703125,-0.1484375,-0.1015625,-0.0078125,0,-0.015625,-0.0625,-0.015625,-0.1015625,-0.1328125,-0.0390625,0.0546875,-0.0703125,-0.0625,0.015625,0.09375,-0.0859375,-0.0703125,-0.0859375,0.1328125,0.140625,-0.0078125,0.0546875,0.0546875,0.125,-0.0078125,-0.09375,0.0234375,0.046875,0.046875,-0.0625,-0.109375,0.0078125,-0.0859375,0.0078125,-0.0625,0.03125,0.1015625,-0.1796875,0.1640625,-0.171875,-0.0625,0.0859375,0.0859375,0.1484375,0.046875,-0.0859375,0.046875,-0.0546875,-0.1015625,-0.03125,-0.0703125,0.0078125,0.1171875,-0.0390625,-0.046875,-0.078125,0.2421875,0.015625,0.046875,0,0.1015625,0.1171875,0,-0.0078125,0.0234375,-0.0390625,0,0.0703125,-0.015625,0.0078125,-0.03125,-0.078125,0.109375,-0.09375,0,-0.046875,-0.03125,-0.0078125,-0.1328125,-0.0859375,-0.0390625,0.015625,-0.015625,0.015625,0.0703125,-0.1484375,0.0234375,0.078125,-0.0703125,0.03125,-0.1484375,-0.0078125,0.1015625,-0.0546875,0.0546875,0.078125,-0.109375,0,0.0078125,0.046875,0.0546875,-0.078125,0,-0.0078125,0.0546875,0.015625,-0.0234375,0.03125,0.0078125,-0.015625,0,-0.0234375,-0.015625,0.03125,0.15625,-0.03125,-0.046875,0.0234375,-0.0234375,0.0234375,0.0078125,0,0.0234375,-0.0234375,0.0390625,-0.046875,-0.109375,-0.015625,0.0390625,0.09375,-0.0234375,-0.03125,0.0078125,0.015625,-0.015625,0.0859375,0.03125,0.0078125,-0.03125,0.0078125,0,0.0546875,-0.0078125,0.078125,-0.03125,0.203125,0.0234375,0.1015625,0.0078125,-0.0078125,0.0546875,-0.015625,0,0,-0.0234375,-0.0390625,-0.078125,-0.0078125,-0.078125,0.0859375,0,-0.015625,0.0078125,-0.0703125,0.0234375,0.015625,-0.0234375,-0.015625,-0.0078125,0,-0.0078125,-0.0390625,0.0078125,-0.015625,0.015625,-0.078125,-0.046875,-0.09375,-0.015625,-0.015625,-0.0390625,-0.03125,-0.046875,0.046875,0.0078125,-0.0859375,0,-0.0859375,0.0546875,-0.0390625,0.015625,0.0078125,-0.03125,-0.0859375,-0.109375,-0.0078125,0.0078125,0.0078125,-0.0078125,-0.03125,0.0234375,-0.0078125,0.0078125,-0.015625,0.09375,-0.03125,-0.015625,-0.0078125,-0.0546875,0,-0.0078125,0.0625,-0.109375,-0.0078125,0.078125,-0.0078125,-0.0234375,-0.015625,0.15625,0.09375,0.1328125,-0.0234375,-0.0546875,-0.0390625,0,0.0234375,-0.0390625,-0.015625,-0.015625,-0.046875,0.046875,0.0390625,-0.0859375,0,0.03125,-0.078125,0.046875,-0.0234375,-0.03125,0.0625,0.046875,0.1171875,0.0078125,0.0546875,-0.0625,-0.03125,0.0703125,0,0.078125,-0.078125,0,0.0390625,0.03125,-0.0703125,0.015625,-0.0546875,-0.015625,-0.0390625,-0.03125,0.078125,0.03125,-0.0546875,0.0234375,0.0625,-0.046875,-0.0234375,-0.0703125,0.1015625,0.0078125,0.046875,0,-0.0390625,0,-0.0078125,-0.0390625,-0.0390625,0,0.03125,0.078125,-0.0234375,0.03125,0.125,0.0078125,0.0078125,0.046875,-0.0234375,-0.046875,0.0234375,-0.0703125,0,0.015625,-0.0078125,-0.09375,-0.09375,0.03125,0.125,-0.015625,0.0546875,-0.0546875,0,-0.0703125,0.015625,0.046875,0.0078125,-0.03125,0.0078125,-0.0703125,-0.0625,-0.0234375,0.046875,-0.0546875,-0.0390625,0.0390625,-0.046875,-0.078125,0.0390625,-0.0078125,0,-0.0078125,0,0.0078125,0.015625,0.0625,-0.09375,0.046875,0.0390625,-0.0546875,0,-0.015625,-0.0078125,0.0078125,-0.078125,0.0703125,0.03125,-0.0546875,-0.0859375,0.0703125,-0.15625,-0.0546875,0.1015625,0,-0.03125,-0.1015625,-0.046875,0.0234375,-0.03125,0.0390625,0.046875,0.0078125,-0.0859375,-0.03125,-0.0625,-0.0078125,-0.0390625,0.0234375,-0.0078125,-0.0078125,-0.046875,-0.0390625,-0.03125,-0.0078125,-0.015625,0.0234375,0.015625,0,0,0.015625,-0.015625,0.0078125,0.0390625,-0.0546875,0,0,-0.0390625,0.0859375,0.015625,0,0.0078125,0.0234375,-0.0390625,-0.015625,-0.0234375,-0.0078125,-0.0234375,-0.0078125,-0.0078125,0,0.03125,-0.015625,-0.015625,0.015625,-0.0390625,0,0.0078125,-0.015625,-0.015625,0.03125,0.0859375,-0.0703125,0.0390625,0.09375,0.0390625,0.03125,0.0859375,-0.0390625,0.09375,-0.015625,0.03125,0.0390625,-0.0234375,0.03125,0.0078125,0.0390625,-0.015625,-0.0234375,0.015625,-0.0078125,0.0546875,-0.0078125,0.015625,-0.03125,0.0546875,0.0234375,-0.0078125,-0.0078125,0.046875,0.0078125,-0.0390625,0,0.03125,-0.0234375,0.0234375,0,0,-0.0234375,0.015625,0.0078125,-0.015625,-0.0078125,0.015625,0.0703125,-0.1328125,0.015625,-0.0546875,-0.015625,-0.0546875,0.0390625,0,-0.015625,0.015625,-0.0390625,0.015625,0.015625,0.015625,-0.0078125,0,-0.0234375,0.078125,0,0.0859375,0.0546875,-0.03125,-0.0078125,-0.0234375,0.0703125,-0.0390625,-0.0546875,-0.0078125,-0.0625,-0.0078125,-0.0234375,-0.0078125,0.015625,-0.0234375,0,-0.0703125,0.015625,-0.03125,-0.109375,0.0234375,0.0078125,-0.015625,0,0,0,0.0859375,0.0078125,-0.046875,-0.0234375,-0.03125,-0.0625,0.09375,0.0703125,-0.0078125,-0.046875,-0.0390625,-0.0234375,0.046875,-0.0078125,0,0.015625,-0.0625,-0.078125,-0.03125,-0.046875,-0.0078125,0.015625,0.0234375,0,0,-0.046875,0,0.046875,0.0234375,-0.0625,0.0078125,-0.0390625,-0.109375,-0.0546875,0,-0.0703125,0.0625,0.0703125,0.0390625,-0.0390625,-0.0625,0.03125,0.0234375,0.0625,0,0.03125,-0.0234375,0,0,-0.0390625,-0.015625,0.0546875,0.03125,0.140625,0.0078125,0,0.015625,0.0390625,-0.046875,-0.078125,0.03125,0.0234375,0.046875,0.0234375,-0.015625,0,0.0546875,-0.0546875,-0.0390625,-0.0703125,0.015625,0,0.0078125,0.0234375,-0.0078125,0.109375,-0.0078125,0,-0.0859375,-0.0546875,-0.03125,0.0703125,-0.0234375,-0.046875,0,0.015625,0.015625,-0.0390625,0.015625,-0.0078125,-0.0546875,-0.0234375,-0.0234375,0.0234375,0.0234375,0.03125,-0.015625,0.0078125,0.03125,-0.03125,0.015625,-0.015625,0.015625,0.0546875,0,-0.046875,-0.046875,-0.0703125,0.109375,-0.0078125,0.0234375,-0.0703125,-0.03125,0.046875,-0.0625,-0.0390625,0.0390625,0.0546875,-0.0625,-0.046875,0.0390625,-0.0625,-0.0078125,-0.0078125,0,0.0546875,0.0546875,-0.015625,0.1015625,-0.0390625,-0.03125,-0.0078125,0.078125,-0.015625,0,0.03125,-0.0546875,0.0078125,-0.015625,-0.0078125,0,0.0234375,-0.0390625,0,-0.03125,-0.0703125,0.1015625,0.015625,-0.0078125,-0.03125,0.015625,-0.0078125,-0.078125,0.03125,-0.03125,-0.0078125,0,0.03125,0,0,0.0078125,-0.03125,0.046875,-0.0078125,-0.015625,0.0234375,0,0.0078125,0.0703125,-0.09375,0.015625,-0.0390625,0.0625,0.078125,0.03125,0.015625,-0.015625,0.0078125,0.03125,0.0078125,0.0390625,0.0859375,-0.03125,0.0234375,-0.0078125,-0.03125,0.0078125,-0.0234375,-0.046875,0.03125,0.0234375,-0.046875,0.015625,0.015625,0.0234375,-0.0546875,0.03125,-0.015625,-0.0390625,-0.0078125,0.125,-0.0546875,0,-0.078125,-0.03125,-0.0234375,0.0078125,-0.03125,-0.0390625,0.0078125,0.015625,0.0078125,-0.0234375,0.0078125,-0.078125,0.03125,0.09375,0.015625,0.0078125,0,0.015625,0.046875,-0.015625,0.0078125,-0.015625,-0.015625,-0.015625,0.0078125,-0.0078125,-0.0703125,-0.0078125,0.015625,-0.0078125,-0.0234375,-0.0703125,0.0546875,0.015625,0,-0.015625,0.0078125,-0.0078125,-0.03125,-0.0234375,-0.03125,-0.046875,0.0234375,0.0390625,0.0078125,-0.0078125,-0.015625,-0.0546875,0.0078125,0.0234375,0.0625,0.015625,-0.0234375,-0.0546875,0.0390625,0,-0.0234375,-0.0078125,0.0703125,0.046875,-0.0234375,-0.0234375,-0.0390625,-0.1328125,0.0625,-0.0078125,0.0390625,0.0078125,-0.046875,-0.0390625,0.015625,0.171875,-0.03125,-0.0703125,0.0234375,-0.0703125,-0.078125,0.046875,0.0078125,0.0546875,0.015625,0.09375,0.21875,-0.109375,-0.078125,-0.0703125,-0.0703125,-0.046875,-0.0234375,0.0078125,-0.0078125,-0.0078125,0.046875,0.0625,-0.0625,0.0234375,-0.0703125,0.09375,-0.015625,-0.0234375,-0.046875,-0.1015625,-0.0625,0.1171875,-0.0390625,0,0.046875,-0.0625,0.0078125,0.078125,0.0234375,-0.09375,-0.09375,-0.03125,0.15625,-0.046875,0.046875,0.140625,0.03125,-0.0078125,0.0625,-0.046875,-0.0859375,-0.0078125,0.0625,0.046875,-0.046875,0.0234375,0.0078125,0.0234375,-0.015625,0,-0.0390625,0.21875,-0.0234375,0.0390625,-0.015625,-0.0625,0,-0.0234375,0.03125,-0.0234375,0.0390625,-0.0546875,-0.0234375,0.0859375,-0.09375,0.0546875,-0.046875,0.015625,-0.0078125,-0.109375,-0.0546875,0.0859375,0.0703125,0.203125,-0.0078125,-0.046875,0.1328125,0.125,0.0234375,-0.0546875,-0.0390625,-0.0859375,-0.0234375,0.15625,0.015625,-0.046875,0.0234375,-0.03125,0.0078125,-0.21875,-0.0234375,-0.046875,0,0.125,-0.03125,0.015625,-0.1484375,0.046875,-0.078125,-0.0078125,-0.03125,-0.0390625,-0.0078125,-0.0234375,0.0390625,0.0234375,-0.015625,-0.0234375,-0.0078125,-0.03125,0.1015625,-0.0234375,-0.0078125,-0.0078125,0.0546875,-0.09375,-0.1015625,-0.03125,-0.0234375,0,0.046875,0.125,0.0234375,-0.0859375,0.0546875,0,0.0078125,-0.0546875,-0.0234375,-0.03125,-0.09375,-0.0078125,-0.0234375,0.03125,0.046875,-0.0078125,0.0703125,0.046875,0.0859375,-0.0859375,0.015625,-0.0390625,-0.0859375,-0.0546875,0,-0.0625,0.0703125,-0.0234375,-0.15625,-0.03125,-0.03125,0.015625,-0.0703125,-0.0234375,-0.015625,0,0.09375,-0.015625,0.046875,0.046875,0.015625,-0.03125,0,-0.015625,-0.0078125,-0.03125,0.078125,-0.1171875,-0.03125,0.0859375,-0.0390625,-0.015625,0.140625,0.0390625,0.0078125,0.1015625,0.0078125,0.0078125,0,-0.0234375,-0.015625,0.015625,0,0.03125,0,-0.03125,-0.03125,-0.0390625,-0.046875,0.015625,-0.03125,-0.078125,0.09375,0,-0.0078125,-0.0078125,0.0078125,0.0625,0.0390625,-0.0234375,-0.015625,-0.0625,-0.0859375,-0.1015625,-0.0390625,-0.078125,-0.0078125,-0.078125,0.078125,-0.046875,0.03125,0,0.125,0.046875,-0.0390625,-0.03125,0.0234375,-0.03125,-0.03125,0.0703125,-0.0078125,-0.0390625,-0.015625,0.0078125,0.0078125,0,-0.046875,0.0078125,-0.0078125,-0.0390625,-0.0703125,0.1875,0.0625,-0.03125,-0.125,0.09375,-0.15625,0.0390625,-0.0078125,0.0234375,0.1328125,-0.078125,0.0625,0.0703125,-0.0234375,0.0625,-0.0859375,0.0234375,0.234375,-0.0078125,-0.0234375,-0.140625,0.0078125,0.0546875,-0.1171875,0.0390625,-0.0390625,0.015625,-0.015625,0.03125,0.1484375,-0.125,0.078125,-0.1171875,0.046875,0.015625,0.3046875,0.125,0.171875,0.1328125,-0.109375,-0.03125,-0.09375,0.015625,0.015625,0.015625,-0.0234375,0.046875,-0.015625,0.0703125,-0.09375,-0.0390625,0.140625,0.03125,0.09375,0.1796875,0.0546875,-0.0546875,-0.0703125,-0.078125,0.03125,0.0078125,-0.125,0.0234375,0,0.03125,0.046875,0.0390625,0.109375,0.0234375,-0.0390625,-0.140625,0.078125,-0.03125,-0.078125,0.09375,-0.0234375,0,0.0703125,0.0078125,0.140625,0.109375,-0.140625,0,0.0234375,0.21875,0,-0.046875,-0.078125,0.140625,-0.0859375,0.0546875,-0.0625,0.046875,-0.03125,-0.015625,0.0078125,-0.109375,0.0625,-0.015625,-0.0859375,0.09375,-0.09375,0.09375,0.0234375,0,0.03125,0.2109375,0.1015625,-0.078125,0.0546875,-0.109375,0.0390625,-0.1328125,0.046875,-0.09375,0.0390625,0.0625,0.2109375,-0.0234375,0.0078125,0.125,-0.09375,0.125,0.125,0.0390625,0.0390625,-0.015625,-0.046875,-0.03125,0.015625,0.0546875,-0.0546875,0.0546875,0.0078125,-0.03125,0.0625,-0.015625,0.015625,-0.046875,0.0078125,0,-0.046875,-0.09375,-0.0078125,0.0078125,0.0390625,-0.0234375,-0.0078125,0.0234375,-0.0390625,0.0625,0.0390625,-0.046875,0.0078125,-0.046875,0.0234375,0.0078125,-0.0078125,-0.03125,-0.03125,0.03125,-0.0234375,0.0234375,0.0546875,-0.0625,0.0234375,0.015625,0,-0.0859375,-0.0546875,-0.0390625,0.0546875,0.0546875,-0.015625,0.0078125,0.046875,0.015625,0.015625,-0.0546875,-0.015625,0.0078125,0.0390625,-0.0390625,0,0.0859375,-0.046875,-0.0234375,0.015625,0.0390625,-0.015625,0,0.03125,0.0234375,-0.0234375,-0.0234375,-0.0078125,0.03125,0,-0.0625,0.0390625,0.0546875,0,0,-0.0234375,0.0234375,0.0390625,0.0078125,-0.046875,-0.0859375,-0.0234375,-0.0625,-0.0390625,-0.015625,-0.0390625,0,-0.03125,-0.046875,0.0234375,-0.046875,0,0,-0.0078125,0.0078125,0.03125,0,-0.0078125,0.03125,-0.0078125,0.03125,-0.0625,-0.0234375,-0.03125,0.0078125,-0.109375,0,-0.0625,-0.03125,-0.0234375,0.03125,0.0078125,0.0390625,0.0234375,-0.0546875,-0.015625,0.0234375,-0.078125,0.0078125,0,-0.0234375,0.0234375,0.0078125,0,0.046875,0,-0.03125,-0.0078125,0.03125,-0.0703125,-0.0703125,-0.171875,-0.109375,0.1328125,-0.015625,0.0234375,-0.0390625,0.0078125,0.0390625,0.1015625,-0.0390625,-0.109375,0.046875,0.3359375,-0.09375,0.140625,-0.0546875,-0.078125,0.0546875,-0.140625,0.0546875,0.0078125,0.1171875,-0.1015625,-0.046875,-0.078125,0.0078125,-0.0703125,0.0859375,0.125,0.03125,-0.078125,-0.078125,0.1171875,-0.0703125,0,-0.1484375,-0.1328125,0.015625,-0.0234375,0.1015625,0.171875,-0.0546875,-0.046875,0.03125,0.0703125,-0.1015625,0.125,0.09375,-0.0078125,0.0703125,-0.1015625,-0.0546875,-0.0703125,-0.140625,0.03125,0.0078125,0.140625,0.1640625,0.1640625,0.1171875,0.1328125,-0.0859375,0.03125,0.15625,0.0546875,0.03125,-0.0546875,-0.09375,0.046875,-0.0078125,0.015625,-0.0390625,-0.0390625,-0.1171875,-0.046875,-0.03125,0.0703125,-0.09375,-0.1015625,-0.03125,-0.0625,0.0859375,-0.09375,0.078125,-0.140625,0.15625,0.0703125,0.015625,0.0625,0.0703125,0.046875,-0.109375,0.109375,0.0234375,-0.1484375,0.0234375,-0.0078125,0.046875,-0.0859375,0,0.1171875,0.0078125,-0.015625,-0.140625,0.0078125,-0.1015625,0.15625,0.0625,-0.03125,-0.0078125,0.1171875,-0.0078125,-0.09375,0.0078125,-0.0546875,0.1015625,0.25,-0.0546875,0.1171875,0.0234375,-0.0625,0.0703125,-0.0625,0.1328125,0.1328125,-0.0234375,0,0,0,-0.0078125,-0.0078125,0.0078125,-0.0078125,-0.0078125,-0.0234375,-0.0234375,0.015625,-0.0234375,0.015625,-0.046875,-0.015625,-0.015625,0.03125,0,-0.03125,0.0078125,-0.03125,-0.03125,0.015625,-0.015625,-0.03125,0,-0.0078125,-0.015625,-0.0078125,-0.015625,0,-0.015625,0.0078125,0,-0.0234375,-0.0234375,-0.0234375,-0.0234375,-0.0234375,-0.0390625,0.0078125,0.0234375,0,0,0.015625,-0.0234375,0,-0.015625,-0.0625,-0.015625,0.03125,0,-0.03125,0,0,0.0625,-0.0078125,-0.015625,0,0,-0.0078125,-0.015625,-0.0234375,0.0234375,0,0.0234375,0.0078125,-0.0234375,-0.0390625,0,0.0078125,0.0234375,-0.015625,-0.0078125,-0.0078125,-0.0078125,-0.015625,0,0.0234375,0,-0.0078125,0,0.015625,-0.03125,-0.0078125,-0.015625,-0.0234375,0,-0.0390625,-0.015625,-0.0234375,0.015625,0,0,-0.03125,-0.0390625,-0.0078125,0.015625,0.0078125,-0.046875,-0.015625,0.015625,0,-0.0234375,0.0546875,-0.0078125,0.0078125,0,-0.015625,-0.0234375,-0.015625,0.0625,-0.03125,-0.0234375,-0.0234375,-0.0078125,-0.03125,-0.0078125,-0.015625,-0.0234375,-0.015625,0,0.0234375,-0.0234375,-0.015625,0.0078125,0.0390625,0.0078125,-0.0078125,0.015625,0,0.0078125,-0.015625,-0.0078125,0.0078125,-0.0625,0.0390625,-0.0078125,0.0078125,-0.015625,0.0234375,0.0234375,0.03125,0.046875,0.0703125,0.015625,0.0078125,0,-0.0234375,-0.015625,0.0078125,0.015625,-0.0078125,-0.015625,0.03125,0.03125,-0.03125,0.0234375,0.0234375,-0.0234375,0.015625,-0.0234375,0,0.0078125,0.0234375,-0.0078125,-0.0390625,0.0546875,-0.015625,0.0078125,0.0546875,-0.0234375,-0.015625,0.0390625,-0.015625,0.03125,-0.03125,0.0078125,-0.0078125,0.046875,-0.0234375,-0.0234375,-0.046875,-0.0078125,0,-0.0390625,-0.0234375,-0.0234375,-0.03125,0.015625,0.0390625,0.0234375,0.0234375,0.015625,0.0078125,0.0078125,-0.0078125,0,-0.03125,0.0078125,-0.0234375,0,-0.0078125,0.015625,0.0078125,0.015625,-0.046875,-0.0078125,-0.0078125,0.015625,-0.0234375,0.015625,-0.015625,0.0078125,-0.0078125,0,-0.0078125,-0.0078125,0.0390625,0.0078125,-0.0078125,-0.03125,0.0078125,-0.03125,-0.015625,-0.0234375,-0.0234375,-0.015625,0.0234375,0.015625,-0.03125,0.015625,-0.0078125,0.0234375,-0.0390625,-0.0078125,-0.0390625,-0.0078125,-0.0234375,0.015625,-0.0234375,0,0.0078125,-0.03125,-0.0234375,-0.0078125,-0.0078125,0.0078125,0.0234375,0.0546875,0.0234375,0.0078125,0.078125,0,0.0390625,-0.03125,0,0.015625,0,-0.0078125,0,0.015625,-0.015625,-0.0234375,0.015625,-0.0078125,-0.015625,-0.015625,-0.0234375,0.0859375,-0.0234375,0,-0.0546875,-0.015625,0.0078125,0,-0.03125,0,0.015625,0.0625,-0.015625,0.015625,0,0.0078125,0.0078125,-0.0078125,0.03125,0,0.0234375,-0.015625,-0.0390625,0.0234375,0.0625,-0.046875,-0.0546875,0.0859375,0.0390625,0.0546875,0.03125,-0.0078125,0.0078125,0,-0.0546875,-0.0234375,0.0234375,-0.0078125,0,0,-0.0078125,0.03125,-0.0078125,-0.0234375,-0.0078125,-0.015625,0.0390625,-0.0390625,0,0.0234375,-0.03125,0,-0.0234375,-0.0234375,-0.015625,-0.0390625,-0.078125,0,0.0546875,-0.0234375,-0.0234375,0.015625,-0.0078125,-0.0234375,-0.0078125,0.0078125,0.0078125,0.0390625,-0.0078125,-0.015625,0.0234375,-0.0390625,0.0234375,-0.0078125,-0.0078125,0.0078125,-0.078125,0,-0.0078125,0,0.015625,-0.015625,-0.015625,-0.0703125,-0.015625,0,-0.0390625,-0.03125,0,-0.03125,-0.0234375,0,-0.0234375,-0.015625,0.03125,0.0078125,-0.0234375,-0.0078125,-0.015625,-0.015625,0.09375,0.0703125,0.046875,0.0234375,0.0625,0,0.0078125,-0.015625,-0.0234375,0.0078125,-0.0078125,0.0078125,0.03125,-0.0078125,0.03125,0,0.1171875,-0.0078125,0.0703125,-0.046875,-0.0234375,-0.0703125,-0.0390625,-0.046875,-0.0859375,0.109375,-0.0234375,0.1171875,0.0546875,-0.015625,-0.1015625,0,-0.1328125,0,0.015625,-0.078125,-0.0078125,-0.03125,0.1015625,-0.015625,0.0078125,0.015625,0,0.0703125,-0.03125,-0.046875,-0.078125,0.0234375,-0.046875,0.0859375,-0.0703125,0,0.0546875,0.015625,0.0546875,0,0.09375,-0.078125,-0.0078125,0.1953125,-0.0390625,-0.03125,0.125,0.015625,0.0546875,-0.03125,-0.0078125,-0.0390625,0.015625,0.0234375,0.1328125,-0.0078125,-0.0390625,0.015625,0,-0.1015625,0.0078125,0.1015625,-0.078125,-0.015625,-0.078125,-0.1171875,-0.0390625,-0.09375,0.046875,0.2890625,-0.0390625,0.0078125,0.0625,-0.0390625,0,-0.0078125,0.0234375,0.015625,0,0.0390625,-0.03125,-0.0078125,-0.078125,-0.0390625,0.0546875,0.0234375,0.078125,-0.0625,0.0078125,-0.0546875,0.0390625,-0.0625,-0.03125,0.015625,-0.0390625,-0.0078125,-0.0625,0.0234375,0.046875,0,0.0078125,0.015625,0.0546875,0.0703125,-0.046875,-0.046875,0.03125,0.0625,0.0234375,-0.015625,0.0703125,-0.015625,-0.015625,0.03125,0,0.09375,0.03125,0,-0.0390625,-0.078125,0.015625,-0.0625,-0.0078125,-0.015625,0.03125,-0.046875,-0.015625,0.0390625,0.0390625,0.03125,0.015625,0.0234375,0.015625,0.03125,0.015625,-0.015625,0,0.046875,-0.0234375,0.0390625,-0.0234375,0.0625,0.046875,-0.0078125,0.015625,-0.0546875,0,0.0078125,-0.046875,-0.0625,0.0234375,-0.0546875,0.0703125,-0.0078125,0.125,-0.015625,-0.03125,0.1015625,0.0078125,0.0078125,0.0078125,0.0078125,-0.0234375,-0.046875,0.0078125,0.0078125,0,-0.015625,-0.0546875,0.0078125,-0.0625,0.109375,0.1015625,0.03125,0.0234375,-0.0078125,-0.03125,0.0390625,0,0.03125,-0.046875,-0.0078125,-0.046875,-0.03125,-0.03125,-0.046875,-0.0234375,0.0234375,0.0390625,0.0078125,-0.046875,0.0703125,-0.0546875,-0.0703125,0,0.0546875,-0.046875,-0.046875,0.0234375,-0.0390625,0,-0.0078125,-0.0234375,0.0234375,0.0234375,-0.0234375,-0.015625,0.1484375,0.0078125,0,-0.046875,0.0546875,0.0390625,-0.015625,-0.1328125,0.0078125,-0.09375,0.03125,0.1015625,-0.0078125,-0.015625,-0.0390625,-0.046875,-0.03125,-0.0625,-0.0078125,0.0859375,0.109375,0.0703125,-0.0703125,0.0078125,-0.03125,0.015625,-0.046875,0.0859375,-0.0078125,0,-0.015625,-0.015625,0.0234375,0.0546875,-0.0390625,-0.0234375,0.015625,-0.0234375,-0.0390625,-0.0078125,-0.0546875,0.0078125,0,-0.03125,-0.078125,-0.0234375,0.0234375,0,0,-0.0234375,-0.0234375,0.046875,0.3046875,-0.03125,0.0625,-0.0234375,-0.078125,0.015625,-0.109375,0.1015625,-0.09375,-0.0234375,-0.0078125,-0.140625,0.0703125,0.09375,0.0625,0.0234375,0.0703125,0.171875,-0.046875,0.078125,-0.1171875,-0.0625,-0.1015625,-0.03125,-0.0546875,0.0234375,0.015625,-0.046875,-0.0859375,-0.078125,0.078125,0.046875,0.109375,-0.046875,0.1015625,0.046875,-0.109375,0.078125,-0.0078125,0.03125,0.0703125,-0.03125,-0.0078125,0.109375,0.109375,-0.1015625,-0.046875,-0.0390625,-0.03125,0.109375,0.1015625,-0.0390625,0.078125,0.2109375,-0.0234375,-0.046875,0.0234375,-0.0859375,-0.0078125,0.0234375,-0.1015625,0.0234375,-0.0546875,0.109375,0.015625,0.171875,-0.1171875,-0.0234375,0,0.109375,0.109375,0.0234375,-0.078125,0.0546875,0.03125,-0.078125,0.0546875,0.109375,-0.0859375,-0.1171875,-0.015625,-0.109375,-0.015625,-0.15625,-0.1640625,-0.0859375,0.046875,0.09375,-0.078125,-0.015625,0.0625,-0.078125,0.0859375,0,-0.0078125,-0.046875,0.0703125,-0.0390625,-0.0078125,-0.03125,-0.0859375,0,0.03125,-0.0859375,0.0703125,-0.0546875,0.0078125,0.0546875,-0.0234375,0.0078125,0.0234375,0.0234375,-0.0625,0.0703125,0.0625,-0.109375,0.1640625,-0.0234375,-0.0390625,0.015625,0.0859375,0.0859375,0.03125,-0.046875,0,-0.015625,0.1484375,-0.0078125,-0.0546875,-0.0078125,-0.015625,0.0234375,0.0078125,0.0390625,-0.015625,0,-0.078125,-0.0546875,0,0.0859375,0.0078125,0.0703125,0.0546875,0.0703125,-0.109375,-0.078125,0.0390625,-0.046875,0.0234375,0.078125,-0.046875,-0.015625,0.0078125,0.03125,-0.0078125,-0.03125,0.0078125,-0.0390625,0.1484375,0.09375,-0.015625,-0.0390625,0.1796875,-0.015625,0.03125,-0.0859375,-0.015625,0.0625,0.0546875,0.0390625,0.0234375,-0.0390625,-0.0234375,-0.0078125,0.0390625,-0.0703125,0.03125,-0.0546875,-0.015625,0.0078125,0.015625,-0.0078125,-0.0078125,0,0.0390625,0,-0.0234375,0.0625,-0.03125,0,-0.1015625,-0.0078125,0.0546875,0.0859375,0.03125,-0.015625,0.015625,-0.0546875,-0.015625,-0.0390625,-0.1484375,-0.015625,0.0390625,-0.0234375,-0.0625,0.015625,-0.0078125,-0.0703125,0.0859375,0,-0.0078125,0.03125,-0.0234375,0.0703125,-0.1015625,0.0546875,0.0234375,0,0.1171875,0.046875,0,0.015625,-0.0390625,0.046875,0.0234375,-0.0078125,0.0703125,0,0,0.078125,-0.0078125,-0.0546875,0.015625,0.09375,0,-0.0546875,-0.0234375,0,0.0078125,0.0390625,0.140625,-0.0546875,-0.03125,-0.0078125,0,0.09375,0.0078125,-0.109375,-0.0078125,0.09375,-0.046875,-0.0234375,0.046875,-0.0234375,-0.125,0.0703125,0.2421875,0.0078125,-0.109375,-0.0234375,-0.0625,0.09375,-0.09375,0.0703125,-0.078125,0.1171875,-0.0390625,-0.0859375,-0.0703125,-0.0546875,0,-0.1015625,0.015625,0.3359375,-0.0390625,0.0703125,0.0703125,0.171875,0.21875,-0.078125,0.03125,0.28125,-0.0546875,0.0625,-0.21875,-0.03125,0.0546875,-0.0234375,0.0546875,-0.078125,0.0234375,-0.0859375,-0.1328125,0.046875,0.125,-0.0625,-0.125,0.125,0,-0.140625,-0.0234375,-0.0625,-0.171875,-0.046875,0.1640625,0.0859375,0,-0.046875,0.1015625,-0.0390625,-0.1171875,-0.0859375,-0.0234375,-0.0625,0.0859375,0.1015625,-0.0390625,0.09375,-0.1953125,0.25,0.203125,0.0546875,-0.0078125,0.1484375,0.0390625,-0.0390625,0.046875,-0.1015625,-0.0390625,0.0703125,-0.0078125,-0.109375,0.015625,-0.15625,-0.03125,-0.0078125,-0.0625,-0.1015625,0.015625,0.03125,0.1328125,-0.0625,-0.078125,-0.140625,0.0390625,0.0625,-0.015625,-0.0859375,-0.1796875,0.0390625,0.09375,0.0546875,-0.1328125,-0.078125,-0.234375,-0.0234375,-0.1484375,0.1640625,0.09375,0.0078125,0.0234375,-0.09375,-0.046875,-0.109375,-0.03125,0,0,0.046875,0.1484375,0.2265625,-0.0078125,0.0546875,0.2265625,-0.140625,-0.03125,-0.09375,0.0078125,-0.09375,0.09375,-0.03125,0.03125,0.0390625,0.03125,0.0546875,0,0,0.03125,0.0234375,0,0.03125,-0.0625,0.03125,0.078125,0.0390625,-0.0546875,-0.0234375,0.0078125,-0.0546875,0.0078125,-0.0546875,0.0546875,0.0078125,-0.046875,0.0390625,-0.109375,-0.03125,-0.0546875,0.0703125,-0.0234375,-0.0234375,0.0625,-0.0078125,-0.015625,0.109375,0.015625,0.015625,-0.0234375,-0.0390625,-0.0390625,-0.1640625,-0.0546875,0.0078125,0.0078125,-0.0625,0.078125,0.0078125,0.03125,-0.015625,-0.0234375,-0.0546875,-0.0390625,0.0625,-0.0625,0.0390625,0.0078125,-0.03125,0.0703125,0.0703125,-0.09375,-0.0078125,-0.046875,0.0546875,-0.015625,-0.078125,0.1953125,-0.0703125,0.078125,-0.0078125,0.078125,-0.1015625,-0.0078125,-0.0859375,0.03125,-0.0703125,-0.0234375,-0.03125,-0.046875,0,0.0078125,0.1484375,0.0078125,-0.015625,0.015625,-0.109375,0.0078125,0,0.0078125,-0.078125,-0.046875,0.03125,0.015625,0.0234375,-0.0078125,0,-0.015625,0.046875,-0.0234375,-0.109375,0.0078125,0.2109375,-0.03125,0.0703125,-0.0859375,0.0234375,-0.0390625,0.109375,0,-0.0859375,-0.0078125,-0.0546875,-0.0546875,-0.0390625,0.0625,0.0234375,-0.09375,0,-0.0625,-0.078125,-0.0703125,-0.015625,-0.03125,0.0703125,0,-0.0078125,-0.03125,-0.0390625,0.0703125,0.0703125,0.125,0.109375,-0.0546875,0.015625,-0.0390625,0.125,-0.0234375,0.0078125,-0.09375,0,0.0234375,0.125,0,0.0234375,0.078125,-0.09375,0.140625,0.0390625,0,-0.0625,-0.0859375,0.078125,-0.015625,-0.0234375,-0.03125,0.03125,-0.15625,-0.1640625,-0.140625,-0.03125,-0.09375,0,0.09375,-0.0078125,-0.09375,-0.015625,0.109375,0.0625,-0.0390625,-0.1796875,0.0859375,0.0625,0.15625,0.1015625,0.015625,-0.03125,0.15625,0.015625,0.09375,0.1328125,0.0546875,0.0390625,-0.046875,0.0625,0.03125,0.1640625,0,0.1015625,0.0234375,0.015625,-0.1015625,-0.109375,0.078125,0.03125,0.1953125,0.078125,0.0234375,0.1796875,0.0078125,0.109375,-0.0078125,0.0546875,-0.0390625,0.046875,-0.0703125,-0.015625,0.1484375,-0.1171875,0.109375,0.0625,-0.0859375,-0.0859375,-0.015625,0.109375,0.0859375,-0.1015625,0.1171875,-0.1015625,-0.140625,-0.078125,-0.078125,0.0703125,0.015625,-0.0078125,0.015625,0.078125,-0.046875,0.1171875,-0.0078125,-0.1328125,-0.078125,-0.0546875,-0.0703125,0.078125,-0.0234375,-0.0390625,-0.1640625,0.1953125,0.078125,-0.0703125,-0.1328125,-0.078125,-0.0859375,-0.0859375,-0.03125,0.0234375,0.0234375,0.0078125,0.0625,-0.046875,-0.03125,-0.046875,-0.078125,-0.0078125,0.0703125,0.09375,0.0546875,-0.0234375,-0.0078125,0,0.0078125,-0.0546875,0.078125,0.0078125,0.0078125,0.015625,0.015625,-0.03125,0,-0.0703125,0.0078125,0.015625,-0.015625,-0.0390625,0,0.0625,-0.03125,0.09375,0.0234375,0,0.09375,0.0078125,-0.109375,0.0078125,0.0546875,0.015625,-0.0546875,-0.046875,-0.1640625,-0.0078125,-0.015625,0.0234375,0,-0.0234375,0.0625,0.03125,-0.0234375,-0.1015625,-0.015625,0.046875,-0.0703125,-0.0546875,-0.0234375,0.1171875,-0.09375,0.03125,0.0078125,-0.0078125,0.015625,0.0703125,-0.0625,-0.078125,0.015625,0,0.0625,0.015625,0,0.03125,0.109375,0.015625,-0.0390625,-0.0546875,-0.078125,0.0859375,0.046875,-0.0078125,0.0078125,0.0390625,0.015625,0.03125,0.03125,0.0390625,0.0234375,-0.015625,0.0078125,-0.0390625,0.015625,0.078125,-0.140625,0.015625,-0.125,-0.0078125,-0.03125,0.125,-0.015625,-0.0546875,0.015625,-0.078125,0.0234375,-0.0390625,0,0.0078125,0.0703125,-0.015625,0.09375,0.0859375,0.046875,-0.0078125,-0.03125,-0.0390625,-0.0625,0.1015625,0.0703125,-0.0234375,0.015625,-0.046875,0.015625,0.0078125,0.0234375,0.015625,0.1015625,0.0078125,-0.0703125,0.171875,-0.03125,-0.09375,0.03125,0.015625,-0.0234375,-0.015625,-0.0078125,0.0703125,0.0625,-0.03125,0.1171875,-0.0390625,0.03125,-0.1015625,0.0625,0.0390625,0,0.03125,0.0234375,-0.015625,0.0703125,0.109375,-0.0234375,-0.0546875,-0.0078125,-0.0546875,0.1640625,0.1171875,-0.078125,0.1875,0.0234375,-0.0390625,-0.046875,0.046875,-0.0078125,0,0.03125,-0.203125,0.0625,-0.09375,0.0625,0.0546875,0.03125,-0.0078125,-0.03125,-0.0546875,0.0625,0.1640625,-0.1171875,0.0546875,-0.03125,-0.0390625,0.0078125,0.046875,-0.03125,0.2109375,0.1171875,-0.1171875,-0.0234375,0.03125,0.0546875,0.109375,0.046875,-0.1171875,0.1796875,-0.015625,0.0703125,-0.03125,-0.15625,0.1953125,0.046875,0.0859375,0.109375,0.015625,0.171875,-0.0859375,-0.0390625,0,0.0390625,-0.0703125,0,-0.015625,0.0859375,0.1484375,0.0703125,0.1328125,-0.140625,0.078125,0.0234375,0.0625,-0.0546875,-0.015625,0.1640625,-0.0625,0.0390625,-0.140625,-0.0546875,0.0546875,0.0078125,0.0390625,0,0.1171875,-0.0546875,-0.078125,-0.0078125,-0.1015625,-0.0703125,-0.0546875,-0.140625,-0.015625,0.0703125,-0.046875,-0.09375,0.03125,-0.1328125,-0.21875,0.015625,0.0234375,0.109375,0.0703125,0.2578125,0.0234375,0.109375,-0.09375,0.1484375,0.0234375,-0.1171875,0.0078125,-0.0078125,0,-0.03125,-0.09375,0.0390625,-0.0078125,-0.0703125,0,-0.03125,0.0234375,0.0390625,0.0546875,-0.0703125,0.0625,0.046875,-0.0234375,0.0546875,0.0078125,-0.03125,0.015625,-0.0546875,-0.0625,-0.0859375,-0.0625,-0.0625,-0.0546875,-0.1015625,-0.015625,-0.0078125,0.1875,-0.03125,-0.0546875,0.015625,-0.125,-0.0546875,0.03125,-0.0546875,0.0234375,0.0703125,0.0078125,-0.03125,0,-0.0078125,-0.0234375,-0.0625,-0.046875,0.0078125,0.0390625,0,0.046875,0.03125,-0.0390625,-0.03125,-0.1640625,0.046875,0.03125,-0.015625,0.0703125,-0.015625,0.078125,0.09375,-0.1796875,-0.0859375,-0.0390625,0,-0.0546875,-0.0078125,-0.0078125,0.0859375,-0.0390625,0.0546875,-0.0390625,-0.0078125,-0.03125,-0.015625,-0.0234375,0.125,0,-0.0234375,0.0078125,-0.015625,-0.0234375,-0.0859375,0.25,0.109375,0,-0.0078125,0.0546875,-0.0390625,0.0625,0,-0.0625,0.0078125,0.0234375,-0.0078125,0.0546875,-0.0078125,-0.09375,-0.0078125,0,0.0078125,-0.015625,-0.0859375,-0.0390625,-0.0078125,0.0078125,0.03125,0.0078125,-0.046875,-0.0625,-0.0859375,0.0625,-0.0625,0.0234375,0.0546875,-0.0234375,-0.015625,0.046875,0.046875,0.09375,-0.0078125,-0.0390625,0,-0.0078125,0.046875,0.0703125,0,-0.09375,-0.0078125,0.078125,0.078125,0,-0.015625,-0.0234375,0.0078125,0.015625,-0.0703125,-0.03125,-0.0546875,0.015625,0.03125,0.03125,-0.0546875,-0.0390625,0.09375,0.078125,0.0078125,0.0078125,0.0390625,0.0390625,0.0234375,-0.0703125,-0.171875,-0.0078125,-0.0078125,-0.03125,0,0.1328125,-0.03125,0.0859375,-0.109375,-0.0078125,0.1953125,0.0078125,-0.0390625,0.0703125,-0.0234375,-0.0078125,0.0859375,0.0703125,-0.0234375,-0.15625,-0.046875,-0.09375,0.0859375,0.1015625,0.0234375,-0.078125,-0.0234375,0.0546875,0.03125,-0.0703125,0.03125,0.0390625,0.046875,-0.078125,0.0234375,-0.0390625,-0.03125,-0.171875,-0.015625,-0.0234375,-0.1015625,-0.09375,0.03125,0.015625,0.0703125,-0.046875,-0.046875,-0.015625,-0.03125,-0.015625,0.0078125,0.109375,-0.046875,-0.0234375,0.03125,-0.078125,0.015625,-0.0390625,-0.03125,0.2109375,0.0234375,-0.015625,0.0234375,-0.1796875,0.0703125,-0.078125,0.03125,-0.1015625,-0.0859375,0.015625,0.0390625,0.125,-0.09375,-0.0078125,0.0234375,-0.03125,-0.1015625,-0.0234375,0,0.1328125,0.0546875,0.046875,-0.09375,0.0078125,-0.015625,0.0625,0.0390625,0.046875,-0.0546875,-0.09375,0.0234375,-0.0625,0,-0.0546875,-0.09375,0.1796875,-0.0703125,-0.078125,-0.0546875,-0.0703125,-0.046875,0.03125,-0.0234375,-0.1015625,-0.015625,-0.015625,0.125,0.1640625,-0.046875,-0.09375,0.078125,0.1484375,-0.03125,0.0703125,-0.0625,-0.0234375,0,0.015625,0,0,0.078125,-0.0078125,0.0703125,-0.0234375,0,0.0390625,0,0.1171875,-0.03125,0.0703125,-0.0234375,0.0390625,0.0078125,-0.0546875,0.0546875,0.0390625,-0.0625,-0.03125,0,-0.0390625,-0.015625,0.078125,0.0703125,0.1171875,0,0.015625,-0.0078125,0.015625,0.0078125,-0.0078125,0.046875,-0.015625,0.046875,0.0234375,0.0234375,0.109375,0.015625,-0.0703125,0.03125,0.0390625,0.0625,0.0703125,0.03125,0.109375,0,-0.09375,0.0234375,-0.0546875,0,-0.09375,0.0390625,-0.0546875,-0.03125,-0.0390625,0.0234375,0.046875,0.0546875,0.0078125,-0.0234375,-0.0859375,0.0859375,-0.046875,-0.1328125,0.015625,0.015625,-0.0859375,-0.0078125,0.0078125,0.0390625,-0.03125,0.0078125,0.0078125,-0.03125,-0.046875,0.0234375,0.0078125,-0.0390625,0.046875,-0.03125,-0.0703125,0.0234375,0,-0.0078125,-0.046875,0,0.015625,0,0.109375,0,0.0078125,0.0546875,-0.046875,0.0078125,-0.0859375,-0.0625,0.0859375,0.046875,0.0859375,-0.015625,0.0390625,-0.0234375,0.03125,-0.0546875,-0.03125,0.015625,-0.0703125,-0.078125,0.0234375,-0.0546875,-0.03125,-0.046875,-0.0078125,0.078125,-0.046875,0.015625,0,0.0234375,-0.015625,-0.0078125,-0.0234375,0.03125,0.015625,0,-0.0078125,0.0234375,-0.1484375,-0.15625,0.0078125,-0.0234375,-0.0078125,0.1796875,0.0546875,-0.046875,0.015625,-0.1484375,0.125,0.0078125,0.078125,0.015625,0,0.0234375,-0.0546875,0.03125,0.0703125,-0.046875,0.1171875,-0.0234375,0.015625,0.0703125,0.1953125,0.015625,0.03125,-0.0390625,-0.03125,0.09375,-0.0703125,-0.046875,0.1796875,0,-0.125,0.15625,0,0.0546875,0.0390625,-0.1640625,0.203125,0,0.0625,0.046875,-0.1171875,-0.1484375,-0.0390625,-0.125,0.1484375,-0.09375,-0.1484375,-0.046875,-0.0234375,-0.125,-0.0546875,0.0234375,-0.15625,-0.109375,0.2890625,0.046875,0.0703125,-0.0625,0.0390625,-0.21875,0.0078125,-0.09375,0.109375,0.171875,0.2109375,0.0703125,-0.140625,-0.0234375,-0.1015625,0.109375,-0.0859375,-0.0234375,0.046875,0.03125,-0.03125,-0.0078125,0.2265625,0.0859375,-0.015625,0.015625,0,-0.1171875,0.1640625,0.171875,0.1953125,-0.03125,-0.0078125,0.0859375,-0.0078125,0.03125,-0.0078125,0.109375,0.0546875,0,0.125,-0.1015625,-0.03125,0.171875,0,-0.1796875,0.1484375,-0.1015625,-0.125,0.109375,0.015625,0.0625,0.1328125,-0.03125,0.0703125,0.140625,0.03125,0.0625,-0.0703125,-0.125,-0.015625,0,-0.078125,0.1875,0.1171875,0.0078125,-0.1875,0.1796875,-0.109375,-0.1328125,0.03125,0.03125,-0.015625,-0.03125,-0.015625,0,0.0078125,-0.015625,0.109375,-0.0078125,0,-0.0234375,0.0078125,-0.0625,0,0,-0.0234375,-0.03125,-0.0078125,-0.046875,-0.03125,-0.0234375,-0.0390625,-0.0078125,-0.0703125,-0.015625,-0.03125,-0.015625,-0.0234375,-0.0625,-0.0078125,0.015625,-0.0546875,0.015625,0.0859375,-0.078125,0.046875,0.03125,-0.1171875,0.0078125,-0.0234375,-0.046875,0.015625,-0.0546875,0.0390625,-0.03125,-0.0859375,-0.03125,-0.125,0.1328125,-0.0390625,-0.0390625,0.0390625,-0.015625,0.0078125,0.0234375,-0.015625,-0.0703125,0.0703125,0.0078125,-0.015625,0.0234375,0.046875,-0.0703125,0.0390625,0.0546875,0,-0.0859375,-0.0078125,-0.015625,-0.0234375,0.1015625,-0.046875,0,-0.0390625,-0.0546875,-0.03125,-0.0078125,0,0.078125,0.015625,0,-0.03125,-0.078125,0.03125,0,0.015625,-0.046875,-0.03125,-0.0390625,-0.046875,0,0,0.046875,0.0859375,-0.046875,-0.046875,-0.0859375,-0.0859375,-0.0625,-0.015625,-0.0546875,-0.1171875,0.09375,0.1484375,0.0078125,0.0703125,0.0078125,-0.015625,0.015625,-0.015625,0.0390625,0.0390625,0,-0.0078125,-0.0390625,0.015625,-0.0078125,0,-0.015625,-0.046875,-0.0078125,0.0234375,-0.0703125,-0.0234375,0.078125,-0.0078125,-0.0703125,-0.015625,-0.0390625,0.0546875,-0.0625,0.03125,-0.078125,-0.0546875,0.140625,0.046875,0.0078125,0.03125,0.0859375,-0.03125,0.0625,-0.046875,-0.0703125,0.0078125,0.015625,-0.078125,-0.0625,0.015625,-0.0625,-0.0390625,0.0234375,0,0.0703125,-0.046875,0.09375,-0.03125,-0.0703125,-0.1796875,-0.015625,-0.0546875,0.03125,0,0.171875,-0.0546875,-0.0390625,0.1328125,0.015625,0.0078125,0.0859375,0.0625,0.1015625,-0.0625,-0.03125,0.046875,-0.0390625,0.0078125,0.0234375,0.0703125,0.0078125,0.125,-0.015625,0.09375,0.0234375,-0.0625,0.1015625,-0.0859375,-0.109375,0.0390625,0.171875,-0.0625,0.0234375,0.03125,0.0546875,-0.0625,-0.1953125,-0.0703125,0.1015625,0.015625,0,-0.0078125,-0.015625,-0.09375,0.0078125,0.0625,-0.015625,-0.03125,0,0.015625,0.03125,0.015625,0.03125,0.078125,0.0625,0.078125,0,0.1796875,-0.0390625,-0.0625,0.1015625,-0.0703125,-0.046875,0.1171875,0.015625,-0.0546875,-0.015625,0.15625,-0.109375,-0.0234375,-0.046875,0.0546875,-0.0546875,-0.078125,-0.109375,0.0859375,0.0234375,-0.015625,-0.0390625,-0.1015625,0,-0.046875,0.0546875,0.1640625,0.1171875,0.03125,-0.0234375,-0.015625,0.0390625,0,-0.109375,0.0546875,-0.0390625,0,0.0703125,-0.09375,0.015625,0.0234375,0.0234375,0.0078125,0,0.015625,-0.046875,0,0,0.0390625,-0.0390625,0.15625,-0.0234375,0.046875,0.0078125,-0.0234375,0.0078125,0.09375,-0.0625,-0.0859375,0.046875,0.109375,-0.1328125,0.0703125,-0.0390625,-0.0234375,0.0234375,-0.0234375,-0.015625,-0.0390625,-0.03125,-0.0078125,0.015625,0.0546875,-0.0078125,0.015625,-0.0859375,0.078125,-0.0234375,-0.0078125,-0.0625,0.0546875,-0.0703125,-0.0390625,-0.1015625,-0.0703125,0.0078125,0.0390625,0.0078125,-0.0859375,-0.0546875,0.0078125,-0.109375,-0.109375,0,0.0078125,-0.0234375,-0.0546875,0.09375,0.0234375,-0.0859375,0.0078125,0.0078125,-0.015625,0.0546875,-0.03125,-0.015625,0.0078125,0.0546875,-0.1171875,0.03125,-0.0234375,0.0625,-0.0078125,0,0.0625,0.0078125,0,0.0078125,0.015625,0.0234375,0,-0.109375,0.125,0.0234375,0.03125,-0.015625,0.0234375,-0.015625,-0.0390625,0.0546875,-0.015625,-0.015625,0,-0.0625,-0.0078125,0,-0.09375,-0.0703125,0.0703125,-0.1640625,-0.0078125,-0.0234375,0.046875,-0.0390625,0.1953125,0.0078125,0.1640625,0.015625,-0.1484375,-0.0078125,0.0546875,-0.015625,-0.0234375,0.078125,-0.1484375,-0.0390625,0.0234375,0.0703125,-0.015625,0.015625,-0.0234375,0,0.046875,0.0234375,-0.0625,0.0625,-0.0234375,0.03125,-0.03125,-0.0390625,0.0625,0.03125,0,0.0234375,0.1640625,0.171875,0.046875,-0.0390625,-0.0625,0.0703125,-0.03125,-0.0546875,0.0078125,-0.015625,0.046875,0.1640625,0.0234375,0.21875,0.0390625,-0.09375,0.03125,0.1015625,0.0078125,0.046875,-0.0390625,-0.1328125,-0.046875,0.0546875,-0.1328125,-0.09375,0.0234375,0.0859375,-0.0078125,0.015625,-0.0234375,-0.15625,-0.0390625,-0.015625,-0.09375,0.140625,-0.0234375,-0.078125,0.0078125,-0.140625,-0.09375,0.015625,0.0546875,0.078125,0.1328125,0,-0.0234375,-0.015625,0.0625,0.0546875,-0.0390625,0.203125,-0.0546875,-0.1015625,-0.0390625,0.0078125,-0.015625,-0.015625,-0.046875,0.1015625,0.0078125,-0.0078125,-0.0625,0.015625,-0.0078125,-0.015625,-0.015625,-0.09375,-0.0390625,0.046875,-0.0546875,-0.078125,-0.0234375,0.1015625,-0.0625,0,-0.046875,-0.0078125,0.046875,-0.140625,-0.0390625,-0.1015625,0.03125,-0.0078125,0.0234375,0.3046875,-0.0703125,-0.0078125,0.0546875,0.0078125,0.0625,0,0.1484375,-0.03125,-0.1484375,-0.0078125,0.015625,0.0859375,-0.0625,0.0390625,-0.046875,0.0078125,-0.078125,-0.046875,-0.1015625,0.078125,0.0625,-0.125,0.09375,-0.0546875,0.0390625,0.0078125,-0.03125,0.0546875,-0.015625,0.0625,0.078125,0.0234375,0.140625,0,-0.09375,-0.078125,0.015625,0.1171875,0,-0.0234375,0.0078125,-0.046875,-0.015625,0.0078125,-0.0625,-0.0078125,0.0078125,-0.046875,0.0625,0.0703125,-0.0078125,0,-0.0625,0,-0.0078125,-0.109375,-0.09375,-0.0390625,0.03125,0.03125,0.03125,-0.03125,0.0234375,-0.03125,0.0390625,0.0625,-0.015625,0,0.125,-0.015625,-0.0390625,0.015625,-0.0703125,-0.0078125,0.1328125,0,-0.0390625,0.21875,-0.015625,0.21875,0.1328125,0.1171875,0.03125,0.0078125,0.0234375,0,0.0078125,0.015625,0.0625,0,-0.03125,0.15625,-0.0390625,-0.03125,-0.015625,-0.03125,0.09375,0.0078125,-0.078125,0.0703125,0.0078125,-0.0078125,0.03125,-0.03125,-0.0625,0.0546875,0.0546875,0.03125,-0.09375,-0.015625,0.015625,0.03125,0.078125,0,0.1328125,-0.078125,-0.0078125,0.0859375,0,-0.078125,0.0625,0,0.0546875,0.09375,-0.0234375,0.015625,0.015625,0,-0.0078125,-0.015625,-0.0234375,-0.0625,0.0546875,0.1171875,0.0625,0,0.015625,0.0703125,-0.0234375,0.0078125,0,-0.0078125,-0.09375,0.0078125,0,-0.015625,-0.03125,0.0390625,0.0078125,-0.078125,0.03125,0.0703125,-0.0859375,-0.0390625,0.015625,-0.0234375,0.0390625,0.015625,0.015625,-0.046875,0.046875,-0.015625,0.0390625,-0.0078125,0,0.0234375,-0.109375,-0.015625,-0.0390625,-0.0859375,0.03125,0.0234375,0.125,-0.03125,-0.109375,-0.0546875,0.0703125,0.0234375,0.03125,-0.015625,-0.0859375,-0.015625,0.0390625,0.1015625,-0.0625,-0.03125,0.0703125,-0.0625,0.0390625,0.03125,0.046875,-0.1640625,0.046875,-0.0078125,0.03125,0,-0.0625,-0.0546875,0.0625,0.0078125,-0.03125,-0.0234375,-0.046875,0.109375,0.109375,0.0859375,-0.0703125,-0.03125,0.0625,0.0703125,0,0.109375,0.09375,-0.015625,-0.03125,0.1640625,0.0859375,-0.0703125,-0.0703125,-0.0234375,-0.03125,0.0234375,0,0.1171875,-0.03125,-0.1015625,-0.0625,-0.078125,0.078125,-0.0234375,0,0.0234375,0.0234375,0.0546875,-0.0234375,-0.03125,0.0234375,-0.0234375,0.0546875,0.0625,0.0078125,0.0546875,-0.0703125,0.0078125,-0.0234375,-0.0234375,-0.0390625,-0.046875,0.046875,-0.015625,0.0859375,-0.0546875,-0.03125,-0.015625,-0.1015625,-0.0859375,0.0625,-0.015625,-0.15625,-0.1484375,0.015625,0.109375,-0.1171875,-0.015625,0.1796875,-0.0234375,-0.0546875,-0.046875,-0.0078125,-0.0546875,-0.09375,0.0234375,-0.078125,-0.0234375,-0.078125,0.171875,0,-0.0703125,0.015625,-0.0078125,0.0078125,-0.046875,-0.0625,0,0.015625,-0.0703125,-0.0234375,0.09375,0.046875,-0.015625,0.0078125,0.0625,-0.015625,-0.0078125,0.0625,-0.0625,0,0,-0.0703125,-0.0078125,0.0234375,0.046875,0.0703125,0.015625,0.0234375,0.109375,0.0234375,0.0078125,-0.015625,0.0703125,-0.0859375,-0.0390625,0.1328125,-0.140625,-0.0234375,0.03125,0.03125,-0.0390625,-0.0078125,0.03125,0.0078125,0,0.0390625,0.0078125,-0.0390625,-0.015625,-0.0546875,0.046875,0.078125,-0.0703125,0.0078125,0.078125,0.0859375,0.0546875,-0.0625,0,-0.03125,0.03125,-0.03125,-0.0234375,0.0703125,0.0390625,0.03125,-0.0234375,-0.0078125,0.015625,-0.0546875,-0.0234375,0,-0.015625,-0.015625,-0.0234375,0.0078125,0.0234375,0,0.0546875,0,0.0078125,0.015625,0.0546875,0,0.0390625,-0.015625,0.09375,-0.015625,0.0078125,0.015625,0,0.0859375,-0.0390625,-0.015625,-0.03125,-0.015625,-0.09375,0.0078125,0.1796875,-0.0390625,0,0.09375,0.0390625,0.140625,-0.0390625,0.0234375,0,0,-0.078125,0,0.0078125,-0.09375,0.015625,-0.078125,0.0625,-0.0546875,-0.0703125,-0.0703125,-0.03125,-0.015625,0.0234375,-0.03125,0,0.0390625,0.015625,-0.0546875,-0.0703125,0.015625,0.0859375,-0.0390625,0.03125,0.0625,0,-0.0078125,0.0546875,0.03125,0.0078125,0,-0.078125,-0.0078125,-0.015625,0.0859375,-0.1640625,0.03125,0.0234375,0.109375,-0.0546875,0.1484375,0.0078125,0.1328125,0.140625,-0.1015625,-0.0078125,0.0703125,-0.1171875,-0.125,0.09375,-0.0703125,-0.09375,0.1015625,0.0234375,-0.0546875,-0.03125,0.0546875,0.1640625,0.0625,0.1484375,-0.125,-0.0703125,-0.078125,-0.09375,-0.046875,0.078125,-0.015625,-0.046875,0.046875,0,-0.015625,-0.046875,-0.0390625,0.078125,-0.140625,0.0859375,-0.0390625,-0.046875,0.234375,-0.1484375,0.0390625,-0.046875,0.03125,-0.171875,0.0625,-0.109375,0.1640625,0.0546875,-0.0546875,-0.0703125,-0.2109375,0,0.1953125,-0.0625,0.1640625,0.03125,0.015625,0.125,0.1640625,0,0.0078125,0.0625,-0.0546875,0.0234375,0.015625,0.046875,0.109375,0.0234375,-0.09375,-0.0078125,-0.0859375,0.0390625,0.1015625,-0.0703125,-0.015625,0.1015625,0.0703125,0.0859375,-0.0078125,0.0078125,-0.140625,-0.1015625,-0.0546875,-0.0390625,0.03125,0.21875,-0.0703125,-0.0546875,-0.0390625,-0.046875,-0.03125,0.1484375,-0.0703125,0.0625,-0.078125,0,-0.0625,0.09375,-0.0703125,0.0234375,0.109375,-0.015625,0.0625,-0.0234375,0.0390625,-0.109375,0.0390625,0.09375,-0.125,-0.0390625,-0.0390625,-0.015625,-0.09375,-0.03125,0.15625,0.1328125,-0.0078125,0.0859375,-0.109375,0.015625,-0.0546875,-0.140625,-0.09375,0.0390625,-0.046875,-0.0078125,0.0078125,-0.0078125,0,0.0078125,0.046875,0.0390625,0.0390625,0.0390625,-0.03125,0.0859375,-0.0078125,0.015625,0.0390625,-0.0078125,-0.0546875,0.0625,0.1015625,-0.0234375,0.0625,0.0234375,0.03125,-0.0546875,0.0390625,-0.03125,0.0234375,-0.015625,0.0234375,0.0625,-0.0234375,-0.0546875,0.015625,-0.015625,0.0234375,0,-0.1328125,0.0390625,0.1328125,0.03125,0,-0.0234375,-0.046875,-0.0390625,0.0390625,0.015625,0.0625,0.0078125,0.1328125,0.0546875,-0.0546875,0.015625,0,-0.0078125,-0.0234375,-0.078125,0.03125,-0.03125,-0.0625,0.0859375,-0.0546875,-0.015625,0.0625,-0.0546875,0.0703125,-0.0078125,0.015625,0.0625,0.046875,0,-0.015625,-0.03125,0.09375,0,0.015625,0.0703125,0.0078125,0,-0.0703125,0.015625,0.0234375,-0.0546875,-0.09375,0.03125,0.0625,0,-0.1171875,-0.078125,-0.0078125,0.0234375,0.1015625,0.0234375,0,0.078125,-0.0390625,0.078125,-0.09375,0.046875,-0.03125,0.1484375,0,-0.0703125,-0.015625,0.0390625,-0.140625,-0.046875,0.0234375,0.0078125,0.0234375,-0.015625,0.0546875,0,0.0078125,-0.0234375,0.125,0.015625,0.0078125,0,0.0234375,0.046875,0.0546875,0.0078125,-0.0234375,0.046875,0.0078125,0,0.015625,0.1875,0.0078125,-0.046875,0.046875,0,0.0234375,0.0234375,0.1484375,0.125,-0.0390625,0,0.046875,0.015625,0.171875,0.0546875,0.015625,0.140625,-0.046875,0.1875,0.0234375,0.078125,-0.0390625,0.0859375,-0.0390625,-0.09375,-0.0703125,-0.1875,-0.0390625,-0.1953125,0.0625,-0.046875,-0.0703125,-0.0546875,0,0.0078125,-0.0546875,-0.0859375,-0.078125,0.0234375,0.015625,0.0078125,-0.046875,-0.015625,0,-0.03125,-0.15625,-0.0859375,-0.0078125,-0.0390625,-0.0234375,0,-0.0078125,0.09375,-0.078125,0,-0.1171875,-0.0859375,0.0703125,-0.140625,-0.1953125,0.0546875,-0.1015625,0.0703125,-0.09375,0.0859375,0.3125,0.109375,0.1171875,-0.0078125,0.078125,0.0546875,0.0078125,-0.0078125,-0.125,-0.0078125,0.1015625,-0.0703125,-0.0390625,0.0546875,-0.0234375,0.0078125,-0.15625,-0.046875,0.265625,0.0234375,-0.078125,-0.1015625,-0.078125,-0.03125,-0.0859375,0.015625,-0.0625,-0.015625,-0.078125,-0.0625,0.1171875,0.0703125,0.1640625,0.046875,0.15625,0.15625,0.0703125,-0.09375,-0.0234375,0,0.03125,0.03125,0.0625,0.09375,0.015625,0.0234375,0.15625,0.015625,0.0078125,0.0234375,0.203125,0.078125,0.109375,-0.1796875,0.046875,0.0703125,-0.1640625,-0.0234375,0.0703125,0.0390625,0.171875,0.109375,-0.0625,-0.0390625,0.015625,0.0234375,-0.046875,0,0.0078125,0,0.03125,0,-0.046875,-0.015625,0.0234375,0,-0.0390625,0.1015625,-0.0234375,0.0078125,0.046875,-0.03125,-0.0234375,0.0546875,0.0859375,-0.015625,0,-0.0234375,0.1171875,0.0859375,-0.015625,0.0078125,-0.015625,-0.078125,-0.0390625,-0.015625,0.046875,0,-0.0390625,0.0078125,-0.0078125,0,0.0390625,0,0.015625,0.0234375,-0.03125,0.09375,-0.0703125,0.015625,0.0546875,0.0078125,0.109375,0.015625,0.0625,0.046875,-0.0859375,-0.015625,0.0078125,0.078125,-0.0546875,0.1171875,-0.09375,0.046875,0.109375,-0.015625,-0.0234375,-0.046875,0.015625,-0.0390625,-0.0234375,0.0859375,-0.0546875,0.03125,-0.03125,0.015625,0.125,0.0390625,0.015625,0.1171875,0,-0.0234375,0.1015625,0.015625,0.0078125,-0.0859375,0.046875,0.0703125,-0.03125,0,0,0.0546875,-0.0234375,0.0234375,0.03125,0.0234375,0,0.0703125,-0.03125,0.0078125,-0.1015625,0.0859375,-0.09375,0.0390625,-0.0390625,0.0390625,0.109375,0.0234375,0.0390625,-0.0078125,0.0703125,0.0234375,-0.09375,0.0078125,0.0859375,0.0703125,-0.1171875,0.0703125,-0.0390625,0.0546875,0.0625,0.0234375,0.0078125,0.0546875,0.03125,0,0.0625,0.03125,-0.046875,-0.0390625,0.0078125,0.1953125,0.0390625,-0.03125,-0.1328125,-0.109375,0,0.0078125,-0.03125,0.046875,0.0703125,0,-0.0859375,0.0859375,0.2109375,0.015625,0.0546875,-0.0703125,-0.1484375,-0.0703125,-0.0078125,-0.0625,-0.0234375,-0.015625,0.1328125,0.0078125,0.0546875,-0.0078125,0.2734375,-0.0078125,-0.015625,-0.0703125,-0.0078125,-0.0546875,0.0390625,0,0,0.0625,0.1796875,-0.1015625,0.078125,-0.09375,0.0625,0.1640625,-0.0625,-0.0625,-0.0625,-0.109375,-0.0625,0.0234375,0.0078125,0.0078125,0.046875,0.0078125,-0.15625,0.0546875,-0.0546875,-0.0625,-0.078125,-0.0859375,0,-0.125,0.046875,-0.1640625,-0.0234375,-0.125,-0.03125,0.1171875,0.09375,-0.0078125,0.0625,0.0234375,-0.109375,-0.0234375,-0.015625,-0.0546875,-0.0546875,-0.1640625,-0.1015625,0.0546875,0.078125,0.09375,0.078125,0.078125,0.0234375,-0.1796875,0.1015625,0.0078125,0.0546875,-0.0546875,-0.078125,0.1171875,0.0234375,0.0078125,-0.03125,0.0234375,-0.0625,0,-0.0234375,-0.03125,0.078125,0.0625,-0.015625,0.0703125,0.0390625,0.109375,0.03125,0.078125,-0.0390625,-0.03125,0.1015625,-0.109375,0.09375,0.125,0.046875,-0.2109375,0.109375,-0.2109375,0.015625,0.1171875,-0.0703125,0.0546875,-0.1484375,-0.0078125,-0.09375,-0.0390625,0.046875,-0.03125,-0.0078125,0.0078125,0.0546875,-0.0390625,-0.015625,0,0.0078125,-0.0078125,0,0,-0.03125,-0.03125,-0.0625,-0.0078125,0.0078125,-0.0703125,0.015625,-0.0078125,0.0859375,-0.0234375,0.0390625,0.0078125,0.0546875,0.046875,0.0234375,-0.046875,0.0390625,0.046875,-0.03125,0.0078125,0.0234375,0,-0.0390625,0,0.046875,0.0390625,-0.0078125,-0.0234375,-0.078125,0.015625,0.0703125,0,-0.0625,0.0078125,-0.0859375,0,0.015625,0.1171875,0.1640625,0.03125,-0.015625,-0.0625,-0.015625,0.046875,-0.0234375,0,0.078125,0.1484375,0.015625,0.0234375,-0.1015625,0.046875,-0.046875,-0.03125,0,0.1171875,0.0078125,-0.0390625,0.015625,-0.046875,-0.0234375,-0.046875,0.109375,-0.03125,0.1171875,0.0234375,0.0234375,-0.0390625,0.015625,-0.03125,-0.015625,0.0078125,0.03125,0,-0.015625,0.015625,0.015625,0,-0.0390625,0,0,0.0078125,-0.0078125,0.0078125,0.0234375,0.0625,-0.0234375,0.15625,-0.015625,0,0.0859375,0.0234375,0.0078125,0.0390625,0.0625,-0.0234375,-0.0078125,-0.015625,0,-0.015625,-0.0625,-0.015625,0.0390625,0.046875,-0.0234375,-0.0390625,-0.078125,-0.0546875,-0.046875,0.046875,0,0.046875,0.015625,-0.0078125,-0.0390625,0.1015625,0.0078125,-0.0625,0.015625,0.1484375,-0.1640625,-0.1015625,-0.0859375,0.03125,0.109375,-0.078125,0.21875,-0.0625,-0.1015625,0.2109375,-0.015625,-0.0859375,0.0234375,-0.0078125,-0.0625,0.015625,0,-0.1015625,0.1015625,-0.078125,0.125,-0.0859375,-0.03125,-0.03125,-0.1328125,-0.0625,-0.0546875,-0.046875,-0.0625,0.0625,-0.0625,0.0078125,-0.0625,-0.0546875,-0.0078125,0.1171875,0.09375,0.0703125,-0.0546875,-0.046875,0.0390625,-0.0234375,0,0.0234375,-0.0859375,0.015625,-0.046875,-0.0390625,0.1171875,-0.0703125,-0.0390625,-0.0390625,0.015625,0.0546875,0.2109375,0.0859375,-0.0625,-0.1171875,-0.0546875,-0.0625,-0.1953125,-0.078125,0.015625,-0.0625,-0.0859375,0,-0.0703125,-0.078125,0.046875,-0.0625,0.1328125,0.015625,-0.1171875,-0.0078125,-0.0703125,0.09375,-0.0390625,0.03125,0.046875,-0.078125,-0.0703125,0.0390625,0.0546875,0.0625,0.015625,-0.0234375,-0.03125,-0.140625,-0.078125,-0.125,-0.0078125,-0.015625,0.1171875,0.09375,-0.0078125,0.015625,0.09375,0.015625,0.015625,-0.0234375,-0.0859375,-0.09375,0.2421875,0.0234375,-0.046875,-0.0859375,0.0078125,0.0078125,0.046875,-0.078125,0,-0.1484375,0.1640625,-0.1328125,0.0859375,-0.0234375,-0.015625,-0.015625,0.125,-0.03125,-0.0703125,-0.1640625,-0.0625,0.109375,-0.078125,-0.0546875,-0.0390625,0,-0.0234375,0.015625,-0.046875,0.0234375,0.0078125,0.0390625,0.03125,-0.0390625,0.078125,0.0078125,0.03125,0.0234375,-0.0234375,0.0234375,0.015625,0.015625,0.0859375,0.03125,-0.0234375,-0.03125,0.0234375,0.0234375,0.03125,0.0703125,0.0390625,0,0.015625,0.0234375,-0.015625,-0.0390625,-0.0234375,-0.015625,-0.0703125,0,0,0.046875,-0.0078125,-0.0234375,-0.0625,-0.0078125,0,-0.015625,0.0625,-0.03125,0.1171875,-0.03125,0.0703125,0.0703125,-0.03125,0.0546875,-0.0625,-0.015625,0,0,-0.0078125,-0.0390625,0.03125,-0.0546875,-0.015625,-0.0390625,0.0078125,-0.0234375,0.0703125,0.140625,0,-0.0234375,-0.0078125,-0.015625,-0.0078125,0.0234375,-0.0390625,-0.03125,0.015625,0.0078125,0.0703125,0.1015625,-0.03125,0.0078125,0.0390625,-0.0703125,-0.0078125,-0.078125,-0.0390625,-0.015625,-0.0078125,0.015625,0.0234375,0,-0.03125,0.046875,0.03125,0.0078125,-0.0078125,0.0078125,-0.03125,0.09375,0.0078125,-0.03125,0.1953125,0.0546875,0.078125,-0.0390625,0.015625,0.015625,0.0234375,0.0234375,-0.0078125,0.015625,-0.0546875,0.0234375,0.03125,-0.03125,-0.0234375,-0.0234375,0.03125,0.03125,0.046875,0.015625,0.015625,0.046875,-0.0546875,-0.0078125,0.09375,0,0,0.0625,-0.140625,-0.1875,-0.0078125,0.0390625,-0.046875,-0.0078125,-0.0078125,0.0546875,-0.0625,-0.015625,0.09375,0.0390625,-0.203125,0.0625,-0.0078125,-0.0078125,0.0234375,-0.0625,-0.09375,-0.015625,0.0078125,0.0234375,-0.0625,0,0.15625,0.046875,0.0625,0.0390625,0.21875,0.1953125,-0.015625,-0.0859375,0.0390625,0.0234375,0.1484375,0.078125,0.015625,-0.046875,0.0234375,0.1171875,0.0703125,-0.1484375,-0.09375,-0.0859375,0.0546875,-0.03125,-0.0859375,-0.03125,-0.03125,0.015625,0.0078125,-0.0078125,-0.0234375,0,-0.1953125,-0.125,-0.1484375,-0.015625,0.09375,0.0703125,0.0859375,0.0546875,0.046875,-0.1171875,0.09375,-0.1015625,-0.09375,-0.0625,0.015625,0.1015625,0.1484375,0.078125,0.078125,0.0703125,0.03125,-0.0078125,-0.0390625,-0.0703125,0.1171875,-0.1171875,0.1015625,0.0859375,0.125,0.0859375,-0.109375,-0.0625,0.0703125,0.0234375,0.0859375,-0.015625,0.125,0,0.0625,-0.046875,0.0234375,-0.0625,-0.1171875,-0.09375,-0.0703125,0.03125,0.0859375,0.046875,-0.109375,-0.1875,-0.046875,-0.234375,0,0.03125,0.078125,-0.0390625,0.15625,0.203125,0.1328125,0.1171875,-0.1640625,0.0703125,0.015625,-0.140625,0.0625,0.1015625,0.0703125,-0.015625,-0.046875,-0.0703125,0.171875,0.046875,0.015625,-0.0078125,-0.046875};

weight_1x1 = '{-0.015625,0.0390625,-0.0078125,0,0.0078125,-0.0078125,-0.0078125,-0.0546875,-0.0546875,-0.015625,-0.0078125,-0.0234375,-0.0234375,-0.015625,0.015625,0.109375,0,0,0.0078125,-0.0078125,0.015625,0.0078125,0.0234375,-0.0078125,0,-0.046875,-0.046875,-0.0234375,-0.015625,-0.0234375,0.0234375,-0.03125,-0.0546875,0,0.03125,0.046875,-0.0234375,-0.0078125,-0.0234375,-0.0234375,-0.046875,0.0234375,-0.03125,0.0234375,-0.0546875,-0.0234375,-0.0546875,-0.0234375,0.03125,0.0234375,-0.0078125,0,-0.0234375,0.0703125,0.0234375,-0.015625,0.0078125,-0.046875,-0.0234375,0,-0.03125,0.0390625,0.0234375,-0.015625,-0.0546875,0.03125,0.046875,-0.046875,-0.0625,0.0078125,0.0859375,-0.0078125,0.0625,-0.015625,0.171875,0,-0.015625,-0.03125,0.046875,0.171875,-0.015625,-0.0625,0.03125,0.0859375,0.046875,-0.0390625,0.0234375,-0.0234375,-0.03125,0.0234375,-0.0546875,-0.0703125,-0.046875,-0.015625,-0.015625,0.015625,0.0078125,0.0234375,0.1015625,0.0703125,-0.0234375,0.0234375,0.109375,-0.0625,-0.0859375,-0.0703125,-0.046875,-0.046875,-0.046875,0.03125,-0.0546875,0.03125,0,-0.015625,0.03125,0.03125,-0.0390625,-0.03125,0.125,0.0234375,-0.0390625,-0.046875,0.015625,-0.03125,-0.046875,0,0.015625,0.046875,-0.0078125,-0.03125,0,-0.046875,0.109375,-0.03125,0.0703125,-0.078125,0.0703125,0.0078125,-0.078125,0.03125,0.0390625,0.0078125,-0.078125,0.0078125,-0.015625,0,-0.03125,-0.0546875,0.0234375,-0.0625,0.0078125,-0.0546875,-0.0234375,-0.0859375,-0.03125,0.0234375,0.015625,-0.0625,0.0625,-0.078125,-0.0078125,0.015625,-0.09375,-0.046875,0.0625,0.03125,-0.03125,0.0859375,-0.0078125,-0.0703125,0.0234375,0.046875,0.03125,-0.0078125,0.0234375,0.046875,0,0,0.015625,0.03125,0.03125,-0.03125,-0.015625,-0.0703125,0.0625,0.125,0.03125,0.0625,0.0546875,-0.03125,0.0234375,-0.0078125,-0.0078125,-0.015625,0.0390625,-0.03125,-0.03125,-0.0078125,0,0.015625,0.0078125,-0.0234375,-0.0234375,-0.0078125,-0.0234375,0.03125,-0.03125,-0.015625,0.03125,-0.0234375,-0.03125,-0.03125,-0.0234375,0.015625,-0.0078125,-0.03125,0.0078125,0.0390625,0.0078125,-0.0078125,-0.015625,-0.03125,0.0234375,0,-0.015625,0.0078125,-0.0703125,0.046875,-0.015625,0.03125,-0.0078125,-0.0234375,-0.0859375,-0.03125,0.0078125,-0.0703125,-0.0390625,-0.0234375,0.0078125,-0.0625,-0.0078125,0.03125,0.0390625,-0.0234375,0.0234375,0.0234375,0.03125,-0.0234375,-0.0703125,-0.078125,0.1328125,-0.1171875,0.0234375,0.1484375,0.0234375,-0.0078125,-0.0390625,0.046875,-0.078125,0.0625,0.1015625,-0.0234375,-0.0078125,0.03125,0.0546875,-0.046875,0.0390625,-0.0078125,0.015625,-0.03125,0,-0.0078125,0.015625,-0.0234375,0.0234375,-0.015625,-0.03125,-0.0859375,-0.0546875,-0.0078125,0.0390625,0.0703125,-0.1015625,-0.0234375,0.03125,-0.015625,0.046875,-0.0625,-0.046875,0,-0.0234375,-0.0625,-0.0625,0,0.0859375,-0.0390625,-0.015625,-0.015625,0.0390625,-0.0390625,0.0078125,0.0390625,-0.0546875,-0.0234375,0.03125,-0.0078125,0,-0.0390625,0.015625,-0.0078125,0.0390625,-0.0390625,-0.0078125,0.015625,-0.015625,-0.0625,-0.0078125,0,0.0703125,0.046875,-0.015625,0.015625,-0.015625,0.03125,-0.046875,-0.015625,0.0625,0.0078125,0.0703125,0,-0.0078125,0.0078125,-0.015625,-0.0078125,0.03125,-0.0546875,0.0078125,0.03125,0,0.0546875,-0.03125,-0.015625,0.0234375,-0.046875,0.015625,-0.0078125,-0.046875,-0.03125,-0.0078125,-0.015625,-0.0234375,0.0078125,0.046875,0.0234375,-0.015625,-0.015625,0.0546875,-0.0078125,-0.015625,0.015625,0.0390625,-0.03125,0.0078125,-0.015625,0.03125,-0.03125,-0.0390625,-0.0078125,0.0234375,0.0625,-0.0390625,0.015625,-0.03125,0.0234375,0.0078125,-0.078125,0.0703125,0,0,-0.0078125,-0.0078125,-0.0234375,-0.0234375,0.015625,0.0390625,0.0078125,-0.0078125,-0.0546875,-0.0234375,0.0234375,-0.0390625,0,0.03125,0.015625,0.046875,0.0234375,0.015625,0.0546875,0.015625,-0.015625,0.0234375,-0.015625,-0.03125,-0.0234375,0.0078125,0.0078125,0.0234375,0.0390625,-0.03125,0.015625,-0.046875,0.0390625,-0.0078125,-0.0625,-0.0234375,-0.0390625,-0.0078125,-0.0078125,-0.0546875,0.015625,0,-0.03125,0.015625,-0.03125,0.0625,0.015625,0.046875,-0.015625,0.0390625,0.0078125,0,-0.078125,0.0078125,-0.015625,-0.078125,0.015625,-0.046875,0.0078125,-0.0234375,-0.0546875,-0.0234375,-0.0078125,-0.0234375,0.03125,0.046875,-0.015625,-0.0234375,-0.0078125,0.015625,0.0078125,0.015625,0.046875,-0.046875,0,-0.0390625,0.0625,-0.0625,0.0078125,-0.015625,0.0625,-0.0625,0.03125,0.0234375,-0.0625,-0.0390625,-0.078125,-0.0546875,-0.0390625,-0.0625,-0.0078125,-0.0390625,0,-0.046875,0.15625,0,0.0703125,0.03125,0.1171875,-0.0625,0.140625,0,-0.0234375,0.0390625,0.046875,-0.109375,0.03125,-0.0078125,-0.03125,0.1484375,0.046875,-0.046875,-0.0234375,0.0390625,-0.0390625,0.0546875,0.03125,-0.0234375,-0.0234375,0,-0.03125,-0.015625,-0.09375,-0.0234375,-0.1015625,-0.046875,-0.0234375,-0.0390625,0.078125,-0.0078125,0.0078125,0,-0.046875,-0.0703125,-0.0234375,0.0625,0.0703125,-0.0390625,0.015625,-0.0546875,-0.0390625,-0.046875,-0.015625,-0.0390625,0.0234375,0.0390625,0.0625,-0.046875,-0.015625,-0.015625,0.046875,0.0546875,0.015625,-0.046875,0.015625,0.03125,0.046875,0,0.0546875,0.0546875,-0.0078125,-0.0234375,-0.0078125,0.0078125,0,-0.0390625,-0.03125,-0.0546875,-0.0234375,0.015625,0,0.0078125,0.03125,0.0859375,0,-0.0234375,-0.0625,0.0078125,0.015625,-0.0234375,-0.1015625,-0.0390625,-0.03125,0.078125,-0.0234375,0.0703125,-0.0078125,-0.0625,-0.0546875,-0.0078125,0.0859375,-0.0234375,-0.03125,0.078125,0.0390625,0.0234375,-0.03125,-0.0234375,0.0390625,-0.0234375,-0.0390625,-0.046875,-0.0390625,-0.0234375,-0.0546875,0.015625,-0.0390625,-0.03125,-0.046875,-0.046875,0.0234375,-0.03125,-0.0078125,-0.0078125,-0.0390625,0.046875,0,0.015625,0,0.0859375,-0.0546875,-0.046875,-0.0078125,0.015625,0.0078125,-0.0625,0.0078125,0.0390625,0.0703125,-0.015625,-0.015625,0.0703125,0,0.015625,-0.0390625,-0.0625,0,-0.0078125,0,-0.046875,0.03125,-0.03125,0.03125,-0.015625,-0.0546875,-0.015625,0.0390625,-0.0546875,0.109375,0.046875,0,-0.0703125,0,-0.0234375,-0.03125,0.0390625,0.03125,0.0234375,-0.0234375,-0.0078125,-0.0234375,-0.0390625,-0.0234375,0.03125,-0.0390625,0,-0.015625,0.015625,-0.046875,-0.0078125,-0.015625,-0.0078125,-0.015625,0.0078125,-0.0078125,-0.046875,0.03125,-0.0234375,0,-0.0234375,-0.0078125,0.0078125,0.0390625,-0.015625,-0.015625,-0.0390625,0.0234375,0.0234375,-0.015625,0,-0.03125,-0.046875,0.015625,0.0546875,-0.015625,0.0546875,0.09375,-0.0390625,0.03125,-0.015625,0.078125,0.078125,0.03125,0,-0.03125,0,-0.046875,0.078125,-0.046875,0.03125,0.015625,0.046875,-0.0390625,-0.078125,-0.1015625,-0.0234375,-0.1015625,-0.0703125,0.03125,0.046875,0.015625,-0.0078125,0.0546875,-0.015625,-0.0703125,0.0234375,0.03125,0.046875,0.0234375,-0.03125,0.046875,-0.03125,0,0,0.015625,-0.0234375,0.0546875,0.0234375,0.015625,-0.046875,0.0078125,0.0234375,0.0625,-0.0390625,-0.0078125,-0.0390625,0.0546875,-0.0703125,0.0546875,0.046875,0.015625,-0.078125,-0.03125,-0.015625,0.0703125,-0.0390625,0.0078125,0.03125,0,-0.0546875,-0.0390625,0.03125,-0.0234375,-0.015625,0,-0.015625,-0.0390625,0.0546875,0,-0.03125,-0.0546875,0.046875,0.015625,0,0.0390625,0,0.0078125,0.0234375,0.03125,0.015625,-0.03125,-0.015625,0.0390625,0.0078125,-0.0390625,-0.015625,-0.046875,-0.03125,-0.0625,-0.0390625,-0.0234375,-0.015625,-0.03125,-0.0078125,-0.0234375,0,-0.03125,-0.0390625,0.109375,-0.0234375,-0.0234375,-0.0390625,0.0234375,-0.03125,0.0234375,0.03125,0.0625,0.03125,-0.03125,-0.015625,0.03125,-0.046875,-0.0390625,0.03125,-0.0546875,-0.046875,-0.046875,-0.0234375,0.0625,-0.015625,0.03125,-0.015625,-0.015625,-0.0078125,0,0,0.0234375,0.015625,-0.0390625,-0.015625,-0.0390625,0.0078125,-0.015625,-0.03125,-0.0546875,-0.015625,-0.0078125,0.03125,0.015625,-0.0078125,-0.0234375,-0.015625,0.0390625,0.09375,-0.0078125,0.03125,0.0234375,-0.0234375,-0.0078125,-0.0390625,0.015625,0.03125,0.0390625,0.0546875,-0.0390625,0.0703125,-0.0625,0,-0.015625,0.0234375,0,0,0.0859375,-0.0078125,0.015625,-0.0234375,0.0078125,0.0390625,-0.0546875,0.0078125,0.0078125,-0.015625,0,-0.0625,0.0078125,-0.0390625,-0.046875,-0.0703125,-0.0234375,-0.0625,0.046875,0.0390625,0.046875,-0.0703125,-0.015625,-0.0078125,0.0234375,0,-0.046875,-0.03125,-0.0078125,0.0625,0,-0.0703125,-0.03125,0.09375,0.015625,-0.0390625,0.0234375,-0.0546875,0,-0.015625,-0.0078125,-0.03125,-0.0390625,0,0,-0.0546875,-0.0390625,0.046875,-0.0234375,-0.0390625,-0.03125,-0.03125,0.015625,0.0703125,0.015625,0.015625,0.0234375,0.015625,-0.0234375,-0.046875,-0.03125,0,-0.0234375,-0.015625,0.0234375,0.0390625,-0.015625,0.0078125,0.015625,0,0.0078125,-0.0234375,-0.0234375,-0.0390625,0.03125,-0.0078125,0,0.0390625,-0.046875,-0.03125,0.03125,0.0234375,-0.0546875,-0.03125,0.0078125,0.0390625,-0.015625,0.046875,0,-0.0390625,0.03125,0.046875,-0.0234375,0.015625,0.0546875,-0.0078125,0,0.0078125,-0.0390625,-0.0234375,-0.0078125,-0.0390625,-0.0625,0.0390625,0.0390625,-0.015625,0,0,0.0703125,-0.046875,0.0234375,0.0625,0.0390625,0.0078125,-0.0703125,-0.0234375,-0.015625,0.0078125,-0.0234375,-0.0390625,0.0390625,-0.0546875,-0.03125,-0.0234375,-0.0234375,0,-0.0234375,-0.0078125,0.0234375,0.078125,0.0234375,-0.0078125,0.03125,-0.015625,0.015625,0.0078125,-0.0234375,-0.0546875,-0.0546875,-0.0390625,-0.046875,-0.09375,0.0390625,0.0703125,0.015625,0.03125,-0.0703125,0.0625,-0.0234375,0.0703125,0.0078125,-0.0546875,-0.015625,-0.0625,-0.015625,0.1015625,0.015625,0,0.03125,0.0390625,0,0.09375,-0.0625,-0.015625,-0.0625,0.0234375,-0.1015625,0,-0.0234375,-0.0546875,-0.03125,-0.0546875,-0.0546875,-0.0859375,-0.0234375,0.125,0.0859375,-0.0625,-0.015625,0.03125,-0.046875,0.046875,-0.015625,-0.015625,0,0.0078125,-0.0234375,0.046875,-0.03125,-0.046875,0,0,0.0234375,0.0078125,-0.0078125,-0.0234375,0.03125,-0.0234375,0.0390625,-0.0390625,0,0,-0.046875,0,-0.046875,0.0234375,-0.0546875,0.03125,-0.0546875,0.0546875,0.03125,0.078125,-0.0234375,0.0703125,-0.0546875,0.015625,-0.0234375,0.0234375,0.0234375,0.0625,0.0234375,-0.0390625,0.0078125,-0.0625,0.0078125,-0.03125,0.015625,-0.03125,-0.0234375,-0.046875,-0.015625,0.015625,-0.0625,0.0390625,-0.0234375,0.046875,-0.0546875,0.0546875,0.03125,0.046875,-0.015625,0.0390625,-0.046875,0.046875,-0.0703125,0.03125,0.0078125,0.015625,-0.0234375,0.0234375,0.046875,0.0078125,-0.015625,-0.046875,0.0546875,0.0859375,0.0390625,-0.078125,0.0546875,0.015625,0.0546875,-0.03125,0,-0.0234375,0,-0.0625,-0.0078125,0.0625,0.078125,-0.0625,-0.03125,0.1640625,0.09375,-0.0390625,-0.0234375,-0.015625,-0.0859375,-0.03125,-0.0625,0.078125,0.015625,-0.046875,-0.0390625,-0.0234375,-0.0078125,-0.0234375,-0.0234375,0.015625,-0.03125,0.0234375,0,-0.015625,0.0078125,0.015625,-0.0078125,-0.0078125,-0.03125,-0.03125,0,-0.03125,0.0078125,-0.0390625,0.0234375,0.0234375,0,-0.0078125,-0.0234375,-0.0078125,0.0078125,0.0078125,-0.0234375,-0.0703125,-0.015625,0.09375,0.109375,-0.03125,-0.015625,0,-0.046875,-0.1328125,0.0625,-0.046875,-0.015625,-0.078125,-0.015625,-0.1484375,0.0234375,0.046875,0.078125,0.0078125,0.015625,-0.046875,0.1875,0.0625,-0.0390625,0.015625,-0.09375,-0.0390625,-0.0234375,0.0234375,0.03125,0.0546875,0.0234375,-0.046875,0.0078125,0.0625,-0.015625,0,0.0234375,-0.0078125,0.0234375,-0.0390625,-0.046875,0,0.046875,0.0390625,-0.0078125,-0.03125,-0.046875,-0.03125,-0.0234375,0.0078125,-0.046875,-0.0390625,-0.0546875,0,0.0078125,0.015625,0.0390625,-0.0234375,0.046875,0,-0.015625,0.0234375,0.078125,-0.0390625,-0.0390625,-0.0625,0.078125,0.0625,0.03125,0.0078125,0.0546875,-0.0703125,-0.03125,-0.046875,0.0234375,0.0078125,-0.0078125,-0.03125,-0.0234375,-0.0078125,0.0546875,0.046875,-0.015625,0.0625,0.0078125,0.0234375,0.0234375,-0.03125,0,0.078125,-0.140625,-0.0546875,0.046875,-0.0234375,0,0.0546875,-0.0234375,0.03125,0.015625,-0.0625,0.03125,0.0234375,-0.046875,0.09375,0.109375,0.015625,-0.0390625,0.03125,-0.03125,0.0703125,-0.015625,-0.0078125,-0.0234375,0,-0.03125,-0.0234375,-0.0078125,0.015625,-0.046875,-0.0703125,0,-0.046875,0.0234375,0.015625,0.0234375,0.0390625,-0.0546875,-0.0078125,0.03125,0.0078125,0.0625,0.0234375,0.0234375,-0.0703125,-0.0390625,0,-0.0390625,-0.0234375,0.0078125,-0.0390625,0.0078125,0.0234375,0.015625,-0.015625,-0.03125,-0.015625,0.03125,-0.1015625,-0.046875,0.046875,0.1484375,0.015625,-0.03125,-0.0234375,-0.0625,-0.015625,0.0234375,-0.0546875,-0.0078125,-0.03125,0.03125,-0.0390625,0.0234375,-0.015625,-0.015625,0.109375,0.015625,0.078125,-0.015625,0.0234375,0.03125,-0.0234375,-0.015625,0.0390625,-0.0078125,-0.0078125,0.0234375,0.0078125,0.0234375,-0.0703125,-0.015625,-0.0625,-0.0703125,0.0078125,-0.0078125,0,-0.0390625,-0.0390625,-0.0078125,-0.0546875,-0.0390625,-0.046875,0.0234375,-0.015625,-0.0390625,-0.0234375,-0.03125,-0.0625,0.0703125,0.078125,0,0.015625,-0.0234375,0.0234375,0.03125,-0.0234375,0.03125,0.015625,0.0078125,0.03125,-0.0078125,-0.0859375,-0.03125,-0.015625,0.03125,-0.0546875,0.03125,0,0,-0.0625,-0.046875,0.03125,-0.0078125,0.0390625,-0.0234375,0.0234375,0.0390625,-0.0390625,-0.0078125,0.0078125,0.0234375,-0.03125,0,0.0078125,0.0546875,0,0.03125,0.0625,-0.0625,-0.0234375,-0.0546875,-0.03125,-0.0078125,-0.0546875,-0.0078125,-0.0078125,-0.0546875,-0.0390625,0.09375,0.0546875,0.078125,-0.0390625,0.1328125,-0.0625,0.0703125,0.0703125,0.015625,-0.0234375,-0.015625,-0.0390625,0.0234375,-0.0390625,0.03125,-0.0390625,0.03125,-0.0546875,0.015625,0,-0.0625,0.078125,0.015625,-0.0234375,-0.03125,-0.0625,-0.046875,0.0234375,0.0234375,0.0625,-0.0234375,-0.0078125,0.015625,-0.0234375,-0.0390625,-0.046875,-0.09375,-0.0625,-0.0625,0.0703125,-0.015625,-0.0078125,-0.0703125,-0.046875,0.046875,0.046875,0.0390625,-0.0390625,0.015625,0.0078125,-0.0078125,0.0078125,0.046875,-0.015625,-0.0390625,-0.0078125,0.078125,-0.0703125,-0.046875,-0.0703125,-0.0078125,-0.0078125,0.0625,0.015625,-0.015625,-0.03125,-0.0078125,-0.015625,0.0078125,-0.0859375,0.1171875,-0.03125,-0.015625,0.0078125,-0.0625,0.0546875,0.0234375,-0.0078125,0.0546875,0.0390625,0,-0.046875,-0.03125,0.0078125,0,0.0390625,0.0625,-0.0078125,0.0078125,0,0.109375,-0.015625,0.0078125,0.0390625,0.046875,-0.0234375,-0.0703125,-0.0703125,-0.0859375,-0.015625,-0.046875,0.0234375,-0.03125,-0.0625,-0.0390625,0.03125,-0.0234375,0.046875,0,0.09375,-0.0234375,-0.0390625,-0.0234375,-0.03125,0.0859375,-0.046875,-0.046875,0.0390625,0.0625,-0.0234375,0.046875,-0.0546875,-0.0546875,0.03125,0.0234375,-0.0390625,-0.0390625,-0.03125,-0.0234375,-0.03125,0.03125,-0.0234375,-0.046875,0,-0.078125,0.0078125,-0.015625,-0.0078125,0,-0.03125,-0.0078125,-0.0078125,-0.0234375,-0.046875,-0.0390625,0,-0.03125,0.015625,0.015625,0.0390625,0.046875,-0.0078125,0,0.046875,0.046875,-0.0390625,-0.0078125,-0.0234375,0.0390625,0.015625,0.0078125,0.0234375,-0.03125,-0.03125,0.0078125,0.0234375,0.0078125,-0.015625,0.0234375,0.015625,-0.0703125,0.0390625,-0.0234375,-0.0390625,-0.0390625,0.109375,0,0,-0.015625,0.0234375,0,0.03125,0.0703125,-0.015625,0,-0.03125,0.03125,-0.03125,-0.0703125,0.0078125,0.0078125,-0.015625,0.046875,-0.0859375,0.03125,-0.0078125,-0.0390625,-0.015625,-0.0078125,0.015625,0.015625,-0.0234375,-0.0546875,0,0,-0.046875,-0.046875,-0.0546875,0.0390625,-0.0546875,-0.015625,0.0234375,0.046875,0.0078125,-0.015625,0.0234375,-0.0234375,0.078125,0.0390625,-0.046875,0.0546875,0,0.0078125,-0.03125,-0.0390625,0.046875,0.0234375,0.0078125,0.0234375,-0.0390625,0.0234375,-0.015625,0.03125,-0.0234375,-0.03125,0.0546875,0.0234375,-0.0078125,0.0234375,0.0390625,0.03125,0.0078125,-0.046875,-0.015625,-0.03125,-0.0234375,-0.046875,0.03125,0,-0.0078125,0.0234375,-0.03125,0,-0.015625,-0.015625,0,0.046875,-0.0234375,0.0625,-0.0234375,0.0703125,0.015625,0.015625,0.0234375,0.015625,0.015625,-0.046875,-0.046875,0.0078125,0.015625,-0.0625,-0.046875,0,-0.046875,0.015625,-0.0390625,-0.03125,0.0390625,0.0625,-0.015625,0.0234375,-0.0625,-0.0390625,-0.015625,0.015625,-0.03125,-0.0703125,-0.015625,-0.0078125,0.0625,0.0390625,0.0859375,-0.0234375,0.0078125,-0.046875,0.0234375,-0.015625,0,-0.0078125,0.0078125,-0.03125,-0.0234375,-0.03125,0.0234375,0.03125,-0.0234375,-0.03125,0.0078125,0.0625,0.03125,0.015625,-0.0390625,-0.03125,-0.0234375,-0.015625,-0.015625,-0.0234375,0,-0.0078125,0.0078125,-0.0078125,0.015625,0.0234375,0.0078125,0.03125,0.015625,-0.015625,0.0234375,0.0078125,-0.0234375,-0.03125,0.0859375,0.0390625,0.0625,-0.03125,-0.0078125,0.0078125,-0.0390625,-0.015625,-0.015625,-0.0546875,-0.03125,0.03125,-0.015625,-0.0390625,0.015625,-0.015625,0.046875,-0.0234375,-0.03125,-0.015625,-0.015625,-0.0234375,-0.015625,-0.0078125,0.0234375,-0.046875,0,-0.0078125,0,0.015625,-0.0625,-0.0390625,0.0234375,-0.0390625,0.03125,-0.0234375,0.0390625,0.015625,0.0234375,-0.046875,-0.046875,-0.0234375,0.0078125,0.0859375,0.03125,-0.015625,-0.03125,-0.0234375,0.0078125,0.046875,0.0078125,-0.046875,0.03125,-0.046875,-0.0078125,0.078125,0.0078125,-0.0390625,-0.0234375,0.03125,-0.0078125,-0.015625,-0.0234375,-0.03125,-0.0234375,-0.0078125,-0.0703125,-0.03125,-0.0390625,-0.0078125,0.09375,0.03125,0.03125,0.046875,-0.0078125,-0.046875,0.0390625,0.0078125,-0.0078125,-0.0703125,0.078125,-0.015625,-0.09375,-0.0078125,0.015625,-0.03125,0.1328125,-0.0390625,0.0859375,0.1015625,0.0078125,0.0078125,-0.0390625,-0.015625,-0.0859375,0.078125,-0.03125,0.0390625,0.0546875,-0.015625,0.078125,0.03125,0.03125,0.0078125,-0.0390625,0,-0.015625,-0.0390625,0.03125,0.015625,0.03125,-0.0234375,0,0.0078125,-0.0390625,-0.078125,-0.015625,0,-0.0078125,0,0.0234375,0.03125,0.0078125,-0.015625,0,0.0234375,0,-0.046875,0.0546875,-0.015625,-0.0234375,0.0546875,0.03125,-0.0390625,-0.0234375,-0.015625,-0.0234375,-0.0546875,0.03125,0.0234375,-0.03125,0.0234375,-0.0234375,0.015625,0,-0.0390625,-0.0078125,-0.03125,-0.015625,0.046875,-0.0546875,0.0234375,-0.0078125,-0.015625,-0.046875,-0.0234375,0.03125,-0.03125,-0.0234375,-0.046875,-0.03125,0.0234375,0.0234375,-0.0234375,0.0078125,0.0078125,0.0078125,0.0078125,0.0234375,0,0.015625,-0.0078125,0.0234375,0.0546875,-0.015625,-0.015625,-0.0078125,-0.046875,0.0390625,0.0390625,0.0546875,-0.0546875,-0.0546875,-0.03125,-0.015625,-0.0234375,-0.0390625,0.0859375,-0.046875,-0.015625,0.046875,-0.03125,0.015625,-0.0390625,-0.0625,0.1171875,-0.0625,0,0.015625,0.1015625,0.015625,0.03125,-0.0703125,0,-0.015625,-0.0234375,0.0234375,-0.0078125,-0.03125,0.0078125,-0.0625,-0.0234375,-0.1171875,0.0546875,0.015625,-0.0390625,0.1015625,0.078125,0.03125,0.125,0,-0.015625,0.015625,-0.0078125,-0.0625,0.0078125,-0.015625,0.015625,-0.0390625,0.1171875,0,0.0546875,0.03125,-0.0078125,-0.078125,0.046875,0.0234375,0.0234375,-0.0859375,-0.046875,-0.0078125,0.0703125,-0.078125,0.046875,0.0390625,-0.0078125,-0.09375,-0.0234375,0.015625,-0.0859375,-0.0546875,0.078125,0,0.0390625,0,-0.03125,-0.03125,-0.03125,-0.046875,0.0625,0.0078125,-0.015625,-0.078125,-0.0234375,-0.0078125,-0.0078125,0.078125,-0.1171875,0.0078125,0.0078125,0.0625,0.109375,-0.0546875,-0.0625,-0.0546875,-0.015625,0.0703125,-0.03125,-0.046875,0.015625,0.046875,-0.046875,0.015625,-0.0390625,0.03125,-0.0234375,-0.046875,0.015625,0.0703125,-0.03125,-0.03125,0.03125,0.015625,0.0078125,0.0703125,-0.046875,-0.03125,0,0.015625,0,0.015625,-0.015625,-0.0625,0,-0.0078125,-0.078125,-0.046875,-0.0546875,0.0859375,0.0703125,-0.1015625,-0.0546875,0.0625,-0.0546875,0.015625,-0.0234375,-0.0234375,0.0390625,0.015625,0.0234375,-0.0234375,-0.015625,0.0859375,-0.015625,0.0234375,-0.046875,0.0234375,0.03125,0,-0.0078125,-0.046875,0.0078125,-0.03125,0.0390625,0.0078125,0.0390625,0,-0.046875,-0.015625,0.0078125,-0.015625,-0.0390625,-0.0234375,-0.015625,-0.046875,0.0625,0.0234375,-0.03125,0,0.03125,0.0078125,0.0078125,0.046875,0.0078125,-0.0078125,-0.03125,0.015625,0.1015625,-0.0390625,-0.015625,0.015625,-0.0234375,-0.015625,-0.0078125,0.015625,0.03125,0.0234375,0.0625,-0.0625,0.1171875,-0.0703125,0.0234375,-0.0234375,-0.0390625,-0.0390625,-0.09375,0.0546875,-0.0390625,0.0234375,0.0078125,-0.03125,-0.0078125,-0.046875,-0.0234375,0,-0.0078125,0,-0.03125,0,-0.0234375,0.015625,0.0078125,-0.0078125,-0.0078125,0.0390625,0.0390625,0,0.0078125,0.0234375,0.0546875,-0.015625,-0.03125,0.0234375,0.015625,-0.0390625,-0.0390625,-0.0234375,0.046875,-0.015625,-0.015625,0.0078125,-0.0234375,-0.0234375,0.015625,-0.0390625,0,0.0078125,-0.0078125,-0.0234375,0.0859375,-0.0234375,-0.0078125,0.0078125,0.0078125,-0.015625,0.0390625,-0.0234375,0.0234375,-0.0390625,-0.0234375,-0.046875,0.03125,-0.0546875,0,-0.0625,0.0625,-0.0546875,-0.015625,0.015625,-0.0703125,0.046875,0.03125,0.0625,-0.0078125,0.046875,-0.0234375,0,-0.0078125,0.0390625,-0.03125,-0.046875,0.015625,0.0234375,0,-0.015625,0.0390625,0.0078125,0.0546875,-0.046875,-0.0390625,0.0234375,0.0625,0.0078125,0.03125,-0.0078125,-0.046875,-0.046875,-0.0546875,0.0234375,-0.0078125,0.0703125,-0.0625,0.015625,0.0703125,-0.015625,-0.03125,0.015625,0.015625,-0.0078125,0.03125,-0.0390625,-0.015625,-0.0390625,0.109375,-0.0234375,0.046875,0.0390625,0.0234375,0.0234375,0,0.015625,-0.0546875,-0.0234375,-0.0546875,-0.046875,-0.015625,-0.0703125,0.0234375,-0.0234375,-0.0234375,-0.015625,-0.03125,-0.0234375,0.0234375,0.0078125,-0.015625,0.015625,0.0234375,0.0234375,-0.03125,-0.015625,-0.03125,0,0.03125,-0.0390625,-0.0078125,0.0625,-0.03125,0.0234375,0.015625,-0.015625,0.0390625,0.015625,0.0234375,0.015625,0.03125,0.0078125,-0.0078125,-0.03125,0.0546875,0.046875,-0.0234375,-0.046875,-0.0078125,0.0078125,-0.015625,-0.0546875,0.0078125,-0.03125,-0.0078125,0.0234375,-0.0390625,0.046875,-0.0078125,-0.0546875,-0.0078125,-0.0390625,0.1015625,0.0390625,0.0390625,-0.0234375,-0.03125,0,-0.015625,0.0703125,0.0390625,-0.015625,-0.046875,0,-0.0625,-0.0546875,-0.0390625,0.0234375,-0.0859375,-0.0234375,0,-0.0546875,0.0078125,-0.0625,0.0078125,-0.078125,-0.015625,0.0078125,-0.015625,0.0078125,0.078125,-0.03125,0.03125,-0.0546875,-0.0390625,-0.078125,-0.0390625,-0.03125,-0.015625,0.0078125,-0.0078125,-0.0625,-0.0390625,-0.0234375,0.015625,-0.015625,-0.046875,-0.0390625,0.078125,0.1640625,0.0078125,-0.046875,0,-0.0234375,-0.0078125,-0.0703125,0.0234375,0.0390625,0.03125,0.1328125,-0.0078125,-0.0078125,-0.0625,-0.015625,0.03125,0.0078125,0.0390625,-0.0390625,-0.0234375,-0.046875,-0.0078125,0.0078125,-0.015625,-0.03125,-0.0625,0.0390625,0.0234375,-0.0703125,-0.015625,-0.0078125,0.078125,-0.0234375,0.0078125,0.1015625,-0.046875,0.0078125,0.0859375,-0.046875,-0.0625,0.0078125,0.1484375,0.046875,-0.0390625,-0.078125,-0.0546875,0.0234375,0.0234375,-0.046875,-0.046875,0.0546875,0,0.0546875,-0.0234375,0.03125,-0.0234375,0.0859375,0.03125,0.046875,-0.046875,-0.0546875,-0.0859375,0.0234375,0.0859375,0.1484375,-0.0625,0.0078125,0.015625,-0.0390625,-0.03125,-0.1015625,-0.09375,-0.078125,0,0.0078125,0,-0.0546875,-0.0234375,-0.0078125,0.0234375,-0.0390625,0.0234375,-0.0703125,-0.046875,-0.046875,0.0234375,-0.015625,-0.015625,-0.0546875,-0.0078125,0.0390625,-0.03125,0.0625,-0.0625,0.0625,-0.0234375,-0.0625,0.078125,-0.078125,-0.0625,0,0.0390625,0,0.0078125,-0.0625,0.0390625,0.0234375,-0.0078125,-0.0546875,-0.0390625,0.03125,-0.0078125,-0.015625,-0.0078125,-0.03125,0,0.0703125,-0.03125,0.0078125,-0.0078125,-0.0234375,-0.03125,0.0078125,0,0.0078125,0.0078125,-0.0234375,0.046875,-0.015625,-0.0859375,-0.0234375,-0.0390625,-0.0078125,0,0.0390625,0.0859375,-0.0078125,-0.015625,0.0390625,0.0234375,0.0234375,0.0078125,-0.03125,0.0078125,-0.0390625,0,-0.046875,0.0234375,-0.015625,0.046875,-0.0234375,-0.03125,0,0.0078125,0,0,0.03125,0.0625,-0.015625,-0.0234375,-0.03125,-0.015625,-0.0078125,-0.0390625,0,0.046875,0.0546875,-0.0703125,0.046875,-0.046875,-0.03125,-0.015625,-0.0078125,0.0234375,0.015625,-0.015625,0.09375,-0.03125,-0.015625,-0.0234375,0.0078125,-0.015625,0.0078125,0.015625,0.0546875,-0.0078125,0.015625,0,-0.0390625,0.0625,-0.0234375,-0.015625,0.03125,-0.0078125,0,-0.0546875,0.0078125,-0.0703125,-0.03125,0.0234375,-0.015625,-0.0234375,-0.0390625,0.03125,0.046875,-0.03125,-0.0390625,0.03125,0.0390625,0.0078125,0.0234375,-0.0078125,0.140625,-0.0703125,-0.015625,0.0390625,0.015625,0.015625,-0.0078125,-0.0546875,0.1171875,0.0234375,0.1171875,-0.015625,-0.0703125,-0.0625,-0.015625,0.0078125,-0.03125,-0.03125,0.015625,-0.0234375,0.0078125,0.0390625,0.0546875,0.0390625,-0.015625,0.0078125,0.0703125,-0.0390625,-0.0234375,0.0234375,-0.03125,-0.0546875,0.1015625,-0.0234375,-0.03125,-0.0078125,0.0390625,-0.0703125,0.046875,-0.0078125,-0.0703125,0.0078125,0,0.015625,-0.0703125,0.015625,0.0625,-0.0078125,0.0078125,-0.0703125,0.03125,0.03125,0.03125,0,0.03125,0.0078125,0.0234375,-0.0625,0.0390625,0.03125,-0.0390625,-0.0625,0.0234375,-0.0078125,-0.0546875,-0.03125,-0.0390625,-0.0078125,-0.046875,0.0859375,0,-0.03125,0.0078125,0.03125,0.03125,-0.03125,0.03125,-0.0390625,0.0078125,-0.015625,0.046875,0.015625,0.0234375,0,0.0546875,-0.0234375,0.03125,0.0078125,0.0078125,-0.0546875,0.015625,0.015625,0.015625,0.0546875,0.015625,-0.015625,-0.0546875,0,-0.03125,-0.046875,0.0546875,0.0234375,0,-0.03125,-0.015625,-0.0390625,-0.046875,-0.046875,0.0703125,-0.046875,0.03125,0.0234375,-0.0390625,0.0234375,-0.0625,-0.0234375,-0.0234375,-0.046875,0.078125,0,0.03125,-0.0390625,0,-0.0390625,-0.03125,-0.0234375,-0.03125,-0.0390625,0.03125,0.0078125,-0.015625,0.0078125,0,0.03125,0.03125,0.015625,-0.0234375,0.0078125,-0.0234375,0,0.0234375,-0.015625,-0.03125,-0.0390625,-0.015625,0.0234375,-0.0078125,-0.03125,0.046875,-0.0390625,0.03125,-0.0390625,-0.0234375,0.0625,-0.0625,0,0.046875,0.046875,0.0390625,0.0234375,-0.0546875,0.0234375,-0.0234375,-0.046875,0.0625,-0.0234375,-0.0078125,0.0390625,-0.03125,-0.03125,-0.046875,-0.0234375,-0.015625,-0.046875,-0.0234375,-0.015625,0.0078125,-0.0546875,-0.015625,0.09375,0.0625,-0.078125,-0.0234375,0,0.0625,0.0390625,-0.015625,-0.03125,0.0078125,-0.03125,-0.0703125,-0.046875,-0.0390625,-0.0078125,0.0078125,0.03125,-0.0234375,0.015625,-0.03125,0,0.0390625,0,-0.015625,-0.0234375,0.0078125,0.109375,-0.03125,-0.0078125,0.0078125,-0.046875,-0.078125,0.046875,-0.0390625,0.0078125,0.015625,0.0078125,0.0546875,-0.0625,-0.0703125,-0.03125,0.03125,0,-0.0390625,0.0234375,-0.0078125,-0.0703125,0.0234375,0.0234375,-0.0859375,-0.0390625,0,0.0390625,-0.03125,-0.015625,0.1015625,-0.109375,0.078125,0.015625,0.03125,-0.0390625,-0.015625,-0.03125,0.0078125,-0.03125,0.109375,0.015625,0.015625,0.015625,0,-0.0078125,0,0.0234375,-0.0234375,-0.03125,-0.0078125,-0.0546875,0.015625,0.015625,-0.0078125,0,-0.0234375,-0.0234375,0.0390625,0.0390625,0.03125,-0.0546875,0.03125,-0.015625,0.0625,-0.0234375,-0.0625,-0.0390625,0.0234375,-0.0625,-0.0703125,0.046875,0.015625,0.0234375,0.03125,0.03125,0.015625,0,0.015625,-0.0078125,-0.0390625,-0.0234375,-0.0078125,0.078125,-0.0078125,-0.015625,0,-0.0390625,-0.0078125,-0.015625,-0.0234375,-0.0390625,0.015625,-0.0390625,-0.0234375,0.0078125,0,0,-0.046875,0.03125,0.0390625,-0.0625,-0.015625,-0.0390625,-0.03125,0.0859375,-0.0234375,0.0234375,-0.0234375,-0.015625,0.0234375,-0.015625,-0.0546875,0.0625,0.015625,0.0390625,0,-0.015625,-0.0078125,0.0390625,-0.0234375,0.03125,-0.0234375,0.015625,0,0.109375,-0.015625,-0.0078125,0.0078125,0,-0.046875,-0.0546875,0.0078125,-0.0390625,0.03125,-0.0234375,0.03125,-0.015625,-0.015625,-0.0390625,-0.046875,-0.0234375,-0.0078125,-0.015625,0.0078125,-0.03125,0.0078125,-0.0234375,0.0234375,-0.015625,0.0078125,0,-0.0390625,-0.0234375,-0.03125,0.0546875,-0.0234375,0.0078125,-0.0546875,0.0390625,0.0078125,0.0234375,0,0.0546875,-0.078125,0,-0.015625,0.046875,0.015625,0.0390625,-0.0546875,-0.0078125,0.0625,0.125,-0.0234375,-0.0390625,0,-0.0234375,-0.078125,-0.0546875,0.0078125,0.0078125,0.015625,0.0234375,-0.0625,-0.0859375,-0.03125,0.015625,0.0390625,-0.0234375,0.1015625,0.09375,-0.0390625,-0.03125,-0.1015625,0.09375,0.1015625,0.03125,0.09375,0.15625,0.0234375,0.0546875,0.0234375,0.0390625,-0.09375,-0.046875,0.0546875,-0.015625,-0.0703125,-0.0390625,-0.0703125,0.015625,-0.03125,0.0390625,-0.0078125,-0.0234375,-0.0390625,-0.015625,-0.0234375,-0.0390625,0.0625,0.0625,0,0.109375,-0.046875,-0.03125,0.0390625,-0.0859375,0,-0.09375,-0.015625,0.015625,0.0546875,0.0859375,-0.046875,-0.015625,-0.0078125,0,0.1015625,0,0.0078125,0.03125,0.0234375,-0.046875,0.0078125,-0.0546875,0,0.015625,-0.0625,-0.0703125,-0.015625,0.0859375,-0.0390625,-0.015625,0.0078125,0.046875,0.046875,-0.078125,0.0546875,0.0625,0.0390625,0.015625,-0.0546875,-0.015625,0.0078125,-0.046875,0.0390625,0.015625,0,-0.0234375,0.0546875,-0.03125,0.0390625,-0.0546875,0.09375,-0.0390625,0.0546875,-0.0078125,0,-0.015625,-0.0078125,-0.0234375,0.03125,0.046875,-0.0078125,0,-0.09375,0.015625,0.015625,-0.0546875,0.0546875,-0.09375,0,-0.03125,-0.078125,-0.0078125,-0.0234375,-0.0078125,-0.03125,0,-0.03125,-0.03125,-0.03125,-0.03125,-0.0390625,0.0703125,-0.046875,0.0234375,0.015625,0.03125,-0.0234375,0.0234375,0.0234375,-0.0234375,-0.0078125,0.015625,0.0546875,0.0390625,-0.0625,-0.0703125,0.015625,0.015625,-0.0234375,-0.015625,0.0078125,0.0234375,-0.0078125,-0.0546875,0.046875,0.015625,-0.0546875,0.03125,-0.0703125,-0.078125,0.046875,-0.0078125,-0.015625,-0.0859375,0.1015625,0.0859375,-0.0625,-0.015625,0.0234375,0.0625,-0.0703125,-0.0078125,0.03125,0.03125,0.015625,0.0234375,0.0078125,0.09375,-0.0625,0.125,0.0546875,-0.015625,0.0078125,-0.0625,-0.09375,0,-0.0234375,-0.015625,0.0546875,-0.015625,-0.0390625,-0.015625,0,0,0.0625,-0.0703125,0.0234375,-0.015625,0.125,-0.0234375,-0.0078125,-0.046875,0.078125,0.1484375,0.046875,-0.046875,-0.015625,0.171875,0.0546875,0.0078125,0.0546875,-0.0546875,-0.015625,0.03125,-0.0078125,-0.1015625,-0.03125,-0.0703125,-0.046875,-0.015625,-0.015625,0.0234375,-0.0078125,-0.109375,0.1015625,0.0234375,0.03125,-0.0234375,-0.03125,0.0234375,0.015625,-0.015625,0,-0.015625,-0.078125,-0.015625,-0.0234375,-0.015625,-0.0078125,0.0390625,0.0546875,-0.0546875,0.0625,-0.0546875,-0.0078125,-0.046875,-0.03125,-0.03125,0,-0.046875,0.1171875,0.0703125,-0.0078125,-0.015625,-0.046875,0.0078125,-0.03125,0.0078125,-0.015625,-0.046875,0.078125,-0.0546875,0.0625,-0.046875,-0.046875,0,-0.015625,0.015625,0,-0.03125,-0.015625,-0.0078125,-0.03125,-0.109375,0,0,-0.0546875,0.078125,-0.0625,0.140625,0.0234375,0.0390625,-0.0078125,0.0546875,-0.0390625,-0.0078125,-0.03125,0.078125,-0.0078125,0.015625,-0.015625,-0.0234375,-0.109375,0.0234375,-0.1015625,-0.0234375,-0.015625,-0.0234375,-0.0234375,-0.015625,0.015625,0.0234375,0.0390625,0.0546875,0.0703125,-0.0078125,0.03125,0.0234375,0.0625,0.078125,0.0703125,-0.0546875,-0.046875,0.09375,-0.0546875,-0.0625,-0.0078125,-0.0234375,-0.0078125,0.0078125,0.015625,0.0078125,-0.015625,-0.0546875,0.046875,-0.015625,-0.0390625,0.0078125,-0.0390625,0.0625,-0.0234375,-0.046875,0.03125,0.03125,-0.0390625,0.046875,0.03125,-0.03125,-0.046875,0,-0.03125,-0.0078125,0.0703125,0.0234375,-0.0078125,0.0078125,0.0234375,-0.03125,0,0.0234375,0.0625,-0.03125,-0.015625,-0.03125,-0.046875,-0.0078125,-0.0546875,0.0390625,0,0,0.015625,0.078125,-0.03125,0.0546875,-0.0078125,-0.0234375,-0.0390625,-0.0234375,0,-0.0390625,0.0078125,-0.0390625,-0.0546875,-0.046875,0.0625,0.078125,-0.015625,-0.046875,0.046875,-0.0546875,0.0078125,0.015625,0.0703125,-0.0625,0.0234375,0.015625,0.0703125,0.0390625,-0.03125,0.015625,0,0.0390625,0.0390625,0.0234375,-0.0546875,-0.0234375,-0.015625,0.0546875,-0.0625,-0.0078125,-0.0234375,-0.0859375,0.046875,0,0.015625,-0.0234375,0.015625,0.015625,0.03125,-0.0625,0.046875,-0.0546875,0.09375,-0.03125,-0.015625,-0.0625,-0.015625,0,-0.0390625,0.0703125,0,0.0703125,-0.03125,-0.0546875,-0.046875,-0.0546875,-0.0390625,-0.0234375,-0.0078125,0.0078125,0.03125,-0.0078125,-0.0234375,0.0390625,0.0546875,-0.015625,-0.0234375,-0.0234375,0.0390625,-0.0546875,-0.03125,-0.0625,-0.015625,0.1328125,0.015625,0.0078125,0.015625,0.0078125,0,0.0234375,0.1015625,0.0234375,0,-0.0078125,0.0234375,0.0234375,-0.015625,0.0234375,-0.0390625,-0.0234375,0.0078125,0,0,0,-0.0078125,-0.0390625,0.0546875,-0.03125,0.03125,0,-0.0390625,0,0.0078125,-0.0078125,0.078125,0.03125,-0.0390625,0.0234375,-0.078125,0.0078125,0.1015625,0.0078125,-0.0546875,0.0703125,-0.0234375,-0.0390625,-0.015625,0,-0.0234375,0.046875,0.0390625,0.0859375,-0.0390625,-0.015625,-0.03125,0.03125,0.0078125,-0.0078125,-0.03125,-0.046875,0.078125,0.1015625,-0.0703125,0.078125,0.0234375,-0.0078125,0.0390625,-0.03125,-0.0625,-0.03125,-0.03125,0.0390625,0.015625,0,-0.015625,0.0703125,0.015625,0.0078125,0.0546875,-0.0234375,0,0.0078125,-0.03125,-0.015625,0.0234375,-0.03125,-0.0078125,0.0390625,-0.0546875,-0.03125,-0.0390625,0.0390625,0.046875,0.0625,-0.0234375,-0.0546875,0.015625,-0.0078125,0,-0.0234375,0.0234375,-0.03125,0.015625,-0.015625,-0.0390625,-0.0234375,0.015625,0.0625,-0.0234375,0.0546875,0,0.0078125,0.0234375,0.046875,-0.0390625,0.0546875,-0.03125,-0.0625,-0.015625,0.0546875,-0.0234375,-0.0234375,-0.0078125,0.0390625,-0.0234375,-0.03125,0.0703125,-0.0703125,-0.015625,0.03125,-0.03125,0.046875,-0.0546875,-0.03125,-0.03125,-0.0625,0.03125,-0.0390625,-0.0390625,0.0703125,0.0703125,0.0234375,0.0234375,0.0703125,0,0.0546875,0.0078125,-0.0546875,0.0078125,-0.03125,-0.03125,0.015625,-0.0703125,-0.0625,-0.0546875,0.1015625,0.0234375,0.0078125,0.078125,0,-0.0546875,-0.0703125,0.03125,-0.015625,0.03125,-0.0078125,0.0078125,-0.03125,0.0234375,0.03125,0.015625,0.015625,-0.046875,0.015625,0.046875,-0.03125,0,0.046875,0,0,-0.0078125,0.03125,-0.0625,0.015625,0.015625,-0.09375,0.0234375,-0.046875,0.0234375,-0.0234375,-0.0390625,0.015625,-0.0078125,0,0.15625,0.015625,0.0078125,-0.0390625,-0.03125,0.1171875,-0.0546875,0.0234375,0.0625,-0.03125,-0.0078125,-0.015625,0.0234375,0.0078125,-0.0078125,-0.0234375,0,-0.0703125,0.03125,0.0078125,0.0546875,0.015625,-0.046875,-0.0234375,0.0625,0.0625,-0.0234375,-0.0546875,-0.0625,0.0234375,0.0625,0,-0.0078125,-0.078125,-0.0390625,0.0234375,-0.0546875,-0.0546875,0.015625,0.0390625,-0.046875,-0.03125,0.125,-0.015625,-0.0703125,0.015625,-0.0625,0.1015625,-0.0703125,-0.0078125,-0.015625,-0.015625,-0.015625,-0.0625,0.0078125,-0.0078125,-0.0390625,0.1171875,0.0546875,-0.0390625,0.0390625,0.015625,-0.0390625,0.0234375,-0.015625,-0.03125,-0.0078125,-0.015625,-0.0234375,0.015625,0.0078125,-0.03125,-0.0078125,-0.0546875,-0.03125,0.03125,0.0390625,-0.03125,0.015625,0.0390625,0.078125,-0.046875,-0.015625,0.0078125,0.0546875,-0.0625,0.03125,0.0234375,-0.0390625,-0.015625,0,-0.0390625,-0.0625,-0.0390625,-0.0234375,-0.03125,-0.0234375,-0.0234375,-0.1015625,0.0234375,0.03125,-0.0546875,0.0703125,0.03125,-0.03125,0.03125,-0.046875,-0.03125,-0.109375,0.0078125,-0.0703125,-0.0390625,0.015625,-0.0390625,-0.0390625,-0.0078125,-0.0078125,0.140625,-0.0625,-0.0625,-0.03125,0.0546875,0.0390625,-0.0859375,-0.0859375,0.0078125,0.015625,-0.078125,0.0234375,-0.0078125,-0.015625,0.015625,-0.0390625,0.03125,0.03125,0.03125,0.0390625,0.0078125,-0.0390625,0,-0.0234375,0.046875,0.015625,0.0078125,-0.0234375,-0.046875,0.0078125,0.03125,0,-0.0078125,-0.03125,0.0078125,-0.03125,-0.015625,0,0.0078125,-0.0234375,-0.0703125,0.03125,-0.015625,0.0078125,-0.0234375,-0.015625,-0.015625,-0.03125,0.015625,-0.015625,0.0078125,-0.046875,0.015625,0,-0.015625,0.03125,-0.015625,0.015625,0.0078125,0,-0.0546875,0.0234375,-0.015625,0.078125,-0.0234375,0.125,0.015625,-0.0703125,-0.0625,-0.078125,0.0234375,-0.015625,-0.0078125,0.0625,0.0703125,0.0234375,0.015625,0.0390625,0.0078125,-0.0078125,0.0078125,-0.046875,0.0234375,-0.0078125,-0.0390625,-0.0078125,0.0390625,-0.0078125,-0.03125,-0.03125,0,-0.015625,-0.015625,-0.0078125,-0.015625,0.0234375,-0.0078125,0.0703125,-0.0546875,0.015625,-0.0390625,0,0,-0.0234375,-0.0625,-0.0703125,-0.0078125,0.09375,0.03125,-0.0390625,-0.0390625,0.0546875,-0.015625,0.09375,-0.0078125,-0.0859375,-0.0234375,-0.0078125,-0.0078125,-0.0234375,0.015625,-0.015625,0.0078125,-0.0390625,0.0234375,0,-0.0234375,-0.015625,0.0234375,0.0234375,0.0234375,-0.0625,0.0234375,-0.0703125,0,0.078125,-0.0390625,0.046875,0.109375,0.0234375,0.078125,0.0234375,0.0234375,-0.0390625,-0.015625,-0.0078125,0.0078125,0.03125,-0.0390625,0.0078125,-0.0234375,0.0078125,0.046875,-0.046875,0.0546875,-0.03125,-0.0390625,0.03125,-0.0078125,-0.0703125,-0.0234375,0.03125,0.03125,0,-0.0703125,-0.0234375,-0.0078125,-0.046875,0.0625,0.0078125,0.0546875,-0.0078125,-0.0078125,-0.046875,-0.0390625,0.03125,0.046875,-0.0390625,0.0234375,-0.046875,-0.015625,0.0234375,0.0234375,-0.0078125,0,-0.0078125,-0.0078125,-0.0078125,0.0625,0.03125,0.0078125,-0.046875,-0.0234375,-0.03125,0.0859375,0,0.0078125,0.0546875,0.03125,-0.0703125,-0.0546875,0.015625,0.0625,-0.0390625,-0.046875,0,0,-0.03125,0.015625,-0.03125,0.015625,-0.015625,0.0078125,-0.03125,-0.03125,0.03125,-0.0078125,-0.0078125,-0.015625,-0.046875,-0.0234375,0.03125,-0.0390625,-0.015625,-0.0078125,0.0546875,0.0234375,-0.0078125,-0.0546875,0,0.03125,-0.015625,0.03125,0.046875,0.03125,0.0078125,-0.015625,-0.0078125,0.015625,-0.046875,-0.0390625,-0.0234375,-0.0078125,-0.03125,-0.015625,-0.0078125,-0.0390625,-0.015625,0.03125,0.0234375,0.0078125,-0.0390625,-0.03125,0.0234375,0.015625,0.03125,0,-0.015625,-0.015625,-0.0234375,-0.0078125,0.03125,0.0390625,-0.0234375,-0.0078125,0.0234375,-0.046875,0.0234375,0.0078125,0.015625,0.015625,0.015625,0,0.0546875,0.0078125,0.0234375,0.078125,-0.0234375,-0.0078125,0.046875,0.015625,-0.015625,-0.0234375,0.03125,0.0078125,0.0390625,-0.0234375,-0.015625,-0.03125,-0.0390625,0.0625,-0.0078125,-0.0625,-0.0078125,-0.0078125,0,-0.0546875,0.015625,-0.0234375,-0.0234375,-0.015625,0,-0.0078125,0,0.03125,-0.03125,-0.015625,0.0390625,-0.0078125,-0.03125,-0.03125,0.03125,0,-0.03125,0.0390625,-0.03125,0.0859375,0.03125,-0.0390625,0.0703125,-0.03125,0.1328125,0.015625,-0.046875,-0.0390625,0.03125,-0.0234375,-0.0390625,-0.0390625,-0.0390625,-0.0390625,-0.046875,0.015625,-0.0078125,0.0078125,-0.0625,0.09375,0.0546875,-0.015625,0.0078125,-0.0234375,0.0546875,-0.046875,0,-0.03125,-0.046875,-0.0390625,-0.0234375,0.0078125,0.0390625,-0.0234375,0.0390625,-0.0078125,-0.046875,-0.046875,-0.0234375,-0.0078125,0.03125,-0.0625,0.015625,-0.03125,-0.0234375,-0.0546875,-0.03125,-0.03125,0.0234375,0.015625,0.0859375,-0.046875,0.046875,-0.015625,0.0703125,0.0859375,-0.015625,-0.0234375,0.03125,-0.0078125,0.015625,0,-0.03125,0.015625,0.0078125,0.0234375,-0.078125,0.046875,-0.046875,-0.0390625,0.0234375,-0.0546875,-0.03125,0,0.0078125,0.0078125,0.0234375,0.0078125,0.078125,-0.0625,-0.0078125,0.0078125,-0.0234375,0.0078125,0.0390625,0.015625,-0.0234375,-0.0078125,-0.0234375,-0.015625,-0.046875,-0.015625,-0.0078125,-0.0078125,-0.015625,-0.046875,0.03125,0.0390625,0.015625,-0.015625,-0.0234375,0.0546875,0.0546875,-0.0234375,-0.03125,-0.046875,0.0625,-0.03125,-0.0234375,0.0703125,0.03125,-0.0234375};

weight_3x3 = '{-0.0234375,0.03125,-0.0078125,-0.0625,-0.0703125,-0.015625,-0.0078125,0.0234375,-0.0234375,-0.0078125,-0.0078125,-0.015625,0,-0.0078125,-0.0078125,0,-0.0078125,-0.0078125,0.0546875,-0.0546875,0.0234375,-0.015625,0.0234375,0.03125,-0.046875,-0.0078125,0.03125,0.0390625,-0.046875,0.046875,-0.0078125,0,0.0625,-0.015625,-0.0390625,-0.0078125,0,-0.0078125,0.0546875,0.015625,-0.0859375,-0.0859375,0,-0.046875,-0.0859375,0.0078125,0.0078125,0,0.0078125,-0.0078125,0.0078125,0.0078125,-0.0078125,-0.0078125,0.078125,-0.03125,0.109375,-0.0546875,-0.015625,0.0078125,-0.0078125,-0.046875,-0.0703125,-0.0625,0,-0.0234375,0.0546875,0.0390625,0.046875,0,-0.046875,-0.03125,0.0078125,-0.09375,0.109375,-0.0234375,-0.1328125,0.09375,0.0078125,-0.046875,-0.0390625,-0.0078125,-0.0390625,0.0078125,-0.0078125,0,0.0390625,-0.0078125,0.03125,0.0234375,0.046875,0.03125,0.0390625,-0.0546875,-0.1015625,0.0078125,0.0546875,0.015625,-0.0390625,-0.0078125,0.0234375,-0.0234375,0,0.0625,0.015625,-0.0234375,-0.03125,-0.03125,-0.015625,0.03125,-0.015625,-0.0234375,0.015625,-0.03125,-0.0078125,0.0234375,0.0078125,-0.0234375,0.046875,0.046875,0.0546875,0.0234375,-0.0390625,0.0078125,-0.0390625,-0.0078125,0,0.09375,0.03125,-0.0234375,0.0078125,0.03125,0,-0.0234375,-0.0234375,-0.015625,0,0,0.078125,0.015625,-0.046875,-0.0078125,0.015625,0.0078125,-0.015625,0.0078125,0,0,0.015625,0.0234375,0,-0.0078125,-0.015625,0,0.0078125,-0.046875,-0.046875,0.0234375,0.0234375,0,-0.0234375,-0.0390625,0.046875,-0.0234375,0.015625,-0.046875,-0.078125,0,-0.03125,-0.046875,-0.0234375,0.046875,-0.03125,-0.015625,0,0.015625,0.03125,-0.046875,-0.0390625,-0.03125,0.0390625,0.0625,0.03125,-0.03125,-0.0078125,-0.015625,0.0546875,-0.0546875,-0.078125,0.0078125,0,-0.03125,0.03125,0.0078125,0.0390625,-0.0078125,-0.0078125,-0.0625,-0.0234375,-0.0234375,0.0546875,-0.015625,-0.015625,0.125,-0.0234375,-0.03125,-0.03125,-0.0078125,-0.0078125,-0.046875,0.015625,-0.0625,0.078125,-0.0078125,0,0.0234375,0.0078125,-0.0546875,0.015625,0.0078125,-0.0390625,0.015625,0.0078125,-0.0546875,-0.0703125,-0.0859375,0,0.09375,-0.0390625,-0.1171875,-0.0703125,0.046875,0.0390625,0.078125,-0.046875,0.03125,-0.078125,-0.0078125,0.0078125,-0.015625,-0.015625,0,-0.0546875,-0.1328125,0.109375,0.0546875,-0.0390625,-0.0078125,-0.0859375,0,0.0078125,0.03125,0.046875,-0.0234375,0.1171875,0.0234375,-0.0703125,-0.078125,0.0390625,0.0078125,-0.0078125,0.03125,0,0.015625,0.0625,-0.078125,-0.1015625,0.0234375,0.0625,0.03125,0.0390625,-0.0078125,0.0546875,-0.0390625,-0.0234375,0,0,0.0078125,-0.0078125,-0.015625,-0.078125,-0.0234375,0.015625,-0.046875,0.0078125,0.0078125,0.0078125,0,0.015625,-0.0078125,0.0078125,-0.03125,-0.0234375,0.015625,0.015625,-0.03125,-0.0546875,-0.015625,0.0078125,0.015625,-0.0078125,0,0.0078125,0.0078125,0.0078125,-0.0078125,-0.0390625,0.0078125,0.0390625,-0.0390625,0.0234375,-0.0703125,-0.0546875,-0.0546875,0,0.0078125,0.0078125,0.0078125,0,-0.0390625,-0.0234375,-0.0078125,-0.015625,-0.046875,-0.0234375,0.0078125,0.0703125,0.015625,-0.0078125,0.015625,-0.0078125,-0.0078125,0.03125,0.0078125,0,-0.0078125,0.0078125,0.0078125,-0.015625,0,0,-0.0078125,-0.015625,-0.0234375,0.0859375,0.015625,-0.015625,0.0703125,0.015625,-0.0625,-0.046875,0.0390625,0.140625,0.1015625,0.0625,0.0078125,0.0234375,-0.0234375,0.046875,-0.0546875,-0.0390625,-0.0078125,-0.0390625,0,-0.03125,-0.0390625,0.046875,-0.0078125,0.0390625,-0.0078125,0.0234375,0,-0.03125,-0.015625,-0.015625,-0.0234375,0,0.0234375,0.0859375,0.0859375,0.0546875,-0.015625,0,-0.0078125,-0.0234375,-0.0703125,-0.046875,0,0.0078125,-0.015625,0.0234375,0.03125,0.0390625,0.0078125,-0.0078125,0.0078125,-0.03125,-0.046875,0.0390625,-0.0078125,0.0078125,-0.015625,0.0234375,-0.0078125,0.015625,0,-0.0078125,-0.0078125,0.015625,-0.0234375,-0.0234375,0.03125,0.1015625,0.0078125,0,0.0078125,0.015625,0.0546875,0,0.0078125,0.0234375,-0.046875,-0.0625,0.0078125,-0.0703125,-0.015625,0.03125,-0.0234375,0.0390625,-0.0078125,-0.0078125,-0.015625,0.0078125,-0.0078125,0.0078125,0,0.0234375,0,0,-0.0078125,-0.0078125,-0.03125,0,-0.046875,-0.0546875,0.0078125,-0.015625,-0.03125,0.0078125,0,-0.0234375,-0.0078125,-0.046875,0.046875,-0.046875,0.0703125,0.046875,-0.015625,0.0078125,0,0.046875,0.03125,0.015625,-0.0390625,-0.0703125,0.0234375,-0.0546875,0.015625,-0.046875,-0.1015625,-0.046875,0.03125,-0.015625,0.0546875,0.0703125,0.03125,0,0.0078125,-0.0546875,0.015625,-0.046875,0.03125,0.0546875,-0.0078125,-0.0703125,-0.0390625,-0.03125,-0.1015625,-0.015625,-0.03125,0.046875,0.0859375,0,-0.046875,0.03125,-0.015625,-0.03125,-0.03125,-0.0078125,-0.0703125,-0.046875,0.0078125,-0.0078125,0.15625,-0.015625,0,-0.0546875,-0.0625,0.0234375,0,-0.0234375,-0.0625,0.03125,-0.03125,-0.0703125,-0.015625,0.046875,0.03125,0.0078125,-0.015625,0.0234375,-0.0078125,0.015625,0.0546875,0.03125,0,-0.0546875,0,-0.0078125,-0.0234375,-0.0625,0.1015625,-0.09375,-0.03125,0.0078125,-0.109375,-0.1015625,0.015625,0.1484375,0.0625,-0.0390625,-0.015625,0.0859375,-0.046875,0.015625,-0.0625,0.0859375,0.0234375,-0.0234375,0.0234375,0.109375,0.0546875,-0.015625,-0.0625,0,-0.0234375,0.015625,-0.0703125,-0.0390625,-0.0546875,-0.0078125,0.0078125,-0.0859375,0.015625,0.0625,-0.015625,-0.0234375,0.03125,-0.0234375,-0.03125,-0.09375,-0.03125,0,-0.015625,0.015625,0.015625,0,-0.0078125,-0.015625,0.09375,0.0078125,0,0.015625,0.046875,-0.0078125,0,-0.0078125,0,0.0078125,-0.0078125,0,0,0.015625,-0.0078125,-0.015625,-0.0078125,-0.0390625,-0.0234375,-0.046875,0.0078125,-0.0234375,0.015625,0.015625,0,-0.03125,0.0234375,0.0234375,-0.0390625,-0.015625,0.0234375,0,0,0.0234375,0.0390625,-0.015625,-0.078125,-0.046875,-0.03125,0,0.03125,-0.0234375,0.0078125,-0.015625,0,0,0,-0.0078125,0.015625,0,-0.0078125,0.0234375,-0.015625,-0.015625,0,-0.0078125,0.0078125,-0.015625,0.0234375,-0.03125,-0.015625,-0.0390625,-0.0390625,0,0.03125,-0.0234375,-0.0234375,-0.0234375,0,-0.0703125,0,0.015625,0,-0.0546875,-0.03125,0.015625,-0.0625,0,0.0078125,-0.0078125,0,0.0234375,0.03125,0.015625,-0.015625,0.0703125,0.015625,-0.0625,0.0078125,0,0.0390625,0.0078125,-0.0078125,-0.0390625,-0.03125,-0.03125,-0.0078125,0.0234375,-0.0078125,0.0234375,-0.0234375,-0.0390625,-0.03125,-0.015625,0.0078125,0.0078125,-0.0078125,-0.0078125,-0.046875,-0.0234375,-0.0078125,0,-0.015625,0,-0.015625,-0.015625,-0.0078125,-0.0234375,0.015625,0,0.078125,-0.0078125,-0.0234375,-0.046875,0.078125,0.0390625,-0.0234375,0.0703125,0.0390625,0.0234375,-0.015625,0.0390625,-0.03125,0,-0.0390625,-0.0859375,-0.015625,-0.015625,0.046875,0.015625,0.015625,0.0078125,-0.015625,0.0078125,-0.015625,-0.015625,-0.0078125,0,0.03125,0.0078125,0.0703125,-0.03125,-0.015625,0.03125,0.0078125,0,-0.03125,0.046875,0,0.015625,0,-0.0078125,0.0234375,0,-0.0234375,-0.03125,0.0234375,-0.015625,-0.0625,0.0546875,0.0234375,-0.0703125,-0.03125,-0.015625,0.0078125,0.0078125,-0.015625,-0.0078125,-0.03125,-0.0546875,-0.03125,-0.03125,-0.0546875,-0.0078125,0.1015625,-0.03125,0.0546875,-0.0234375,-0.0234375,0,-0.0390625,0.0078125,-0.0390625,0.015625,-0.03125,-0.0234375,0.046875,-0.03125,0,-0.03125,-0.046875,0.015625,0.0234375,-0.015625,-0.046875,0,-0.046875,0.046875,0.0234375,-0.0078125,0.0234375,-0.046875,-0.046875,0,0.0078125,-0.0390625,0.046875,0.015625,-0.0234375,-0.0703125,0.0078125,-0.0078125,0.0234375,0.046875,-0.015625,0.140625,-0.0078125,-0.015625,-0.109375,-0.0234375,-0.0234375,0.015625,-0.0625,-0.015625,-0.1015625,-0.03125,-0.0390625,0.0703125,0.078125,-0.0234375,-0.046875,-0.046875,-0.0078125,-0.015625,0.0390625,0.0390625,0.0390625,-0.1484375,-0.015625,0.078125,-0.0078125,0.0234375,0.0078125,-0.046875,0.0078125,0.0078125,-0.0390625,-0.046875,-0.0703125,-0.0234375,-0.015625,0.078125,0,0.0234375,-0.046875,-0.0078125,-0.0234375,-0.03125,0,-0.046875,0.0390625,-0.0546875,-0.03125,-0.0234375,-0.015625,-0.03125,0.03125,0.0078125,-0.0234375,0.140625,-0.0078125,-0.03125,-0.0390625,-0.0234375,-0.0234375,0,0.0546875,0.0234375,-0.0078125,0.0390625,0.015625,0.015625,0.1015625,-0.046875,-0.0078125,-0.0078125,-0.0078125,0.0078125,0.0234375,-0.03125,-0.015625,-0.015625,0.0078125,-0.015625,0.0234375,0,0.0078125,-0.0390625,-0.0625,-0.0234375,-0.015625,-0.015625,-0.0234375,0.0859375,-0.0625,-0.0078125,-0.046875,0.0390625,-0.0078125,-0.0078125,-0.03125,0.0234375,-0.0859375,-0.0546875,-0.0546875,-0.0234375,0.0859375,-0.0703125,0.0078125,0.046875,0.0078125,-0.0078125,-0.0078125,0.0078125,0,-0.015625,-0.0078125,0,-0.015625,-0.03125,0.03125,-0.03125,0.1328125,0.1015625,-0.078125,-0.078125,-0.0546875,-0.0078125,0,0.1328125,-0.015625,-0.0859375,-0.125,0.0390625,0.015625,0.1171875,0.0390625,-0.015625,-0.046875,-0.0390625,-0.03125,0.0234375,0,0.015625,0.140625,0.0390625,-0.015625,-0.0390625,-0.015625,-0.046875,-0.03125,0.015625,0.015625,-0.0390625,-0.0234375,0.046875,0.0390625,-0.0078125,0.0390625,0.015625,0.0390625,-0.0234375,-0.0390625,-0.078125,-0.03125,0.0703125,-0.0234375,-0.03125,0.0703125,0,-0.046875,0.0078125,-0.0390625,-0.015625,0.0078125,0.0859375,-0.03125,-0.015625,0,-0.0234375,0.03125,0.015625,-0.0234375,0,-0.0546875,0.0546875,0.015625,-0.03125,-0.03125,0,-0.0390625,0.0078125,0.03125,-0.0078125,0.0078125,0.1171875,-0.03125,0.0234375,-0.078125,-0.0625,0.0703125,-0.0625,0.0390625,-0.0390625,0,-0.125,0.1015625,-0.0625,0.0703125,0,-0.0078125,-0.0078125,-0.015625,0,-0.015625,0.015625,0,-0.015625,-0.0546875,0.140625,0.046875,0.0078125,0.0234375,0.015625,-0.03125,-0.046875,-0.0234375,-0.015625,0.09375,0.0546875,-0.0390625,-0.0234375,0,-0.0078125,0.03125,-0.0078125,-0.046875,-0.140625,-0.09375,-0.109375,0.0234375,0.015625,0.078125,-0.0234375,-0.046875,-0.0078125,-0.078125,-0.0078125,0,-0.0078125,0.0703125,-0.03125,-0.0234375,-0.015625,-0.0390625,0.0703125,0.015625,-0.1015625,-0.0234375,-0.1171875,-0.0546875,-0.0703125,0.0078125,-0.0390625,0.0078125,-0.03125,-0.0078125,0.03125,0.0234375,-0.0234375,-0.0546875,0.109375,0.015625,0.0546875,-0.0078125,-0.0234375,-0.0234375,-0.0390625,-0.015625,-0.015625,-0.09375,0.0703125,-0.03125,0.015625,0.015625,0.0703125,-0.0546875,-0.015625,-0.109375,-0.125,-0.0078125,-0.1015625,-0.0625,-0.0546875,-0.078125,0.0625,0.0234375,0.0234375,-0.0078125,-0.0234375,-0.0234375,0.0859375,-0.0546875,-0.0234375,0.015625,-0.0234375,0.0546875,-0.0234375,-0.0859375,-0.0234375,-0.0078125,0.0234375,0.0859375,-0.0078125,0.0390625,-0.03125,-0.0078125,-0.0546875,-0.03125,-0.046875,0.03125,-0.0703125,0.0859375,0,0.0078125,-0.0703125,-0.0703125,0.125,-0.03125,0.0234375,-0.140625,0.03125,-0.0390625,-0.125,0.0625,0.0625,0.0234375,0.046875,-0.109375,-0.109375,-0.0703125,0.015625,0.03125,0.0234375,-0.109375,0.1484375,-0.046875,0.0078125,-0.078125,-0.0078125,-0.0546875,0.03125,0.046875,-0.015625,-0.015625,0.0234375,0.0078125,-0.015625,0,0.0390625,0.0703125,0.015625,-0.0078125,0.0078125,-0.0078125,0.015625,-0.0078125,0,-0.0078125,0.0078125,0.0078125,0,0.0078125,-0.0234375,-0.0234375,-0.0078125,-0.0390625,0.0078125,-0.0390625,0.0234375,0,0.0234375,0,0,0.0078125,0.0078125,-0.0234375,-0.046875,0.0078125,0.015625,-0.0078125,-0.0078125,0.0078125,-0.015625,-0.0625,-0.0234375,-0.0546875,0.03125,0.0078125,0,-0.0078125,0.0078125,0,0.0078125,0,0,0,0,-0.0234375,0.0078125,0.015625,-0.0234375,-0.015625,0.0390625,-0.046875,0.0703125,-0.0078125,0.0703125,0.015625,0.015625,0.03125,-0.015625,0,-0.0078125,0.015625,-0.0078125,-0.0390625,-0.0234375,0,-0.0234375,-0.015625,0.015625,0,-0.015625,0.0078125,-0.0078125,-0.0078125,0,0.0078125,0.0078125,-0.015625,-0.0390625,-0.015625,-0.0390625,-0.015625,-0.015625,-0.015625,-0.03125,0.0078125,-0.0234375,0.015625,-0.0234375,0.0078125,-0.0078125,0.0234375,0,-0.015625,-0.0078125,0.015625,0.0078125,-0.0078125,0,0.03125,0.015625,-0.0078125,-0.0234375,0.0078125,0,-0.0078125,0.03125,-0.015625,0.0234375,0,-0.03125,-0.0234375,0,-0.0078125,0.03125,-0.0078125,-0.03125,0.015625,0.0078125,-0.0234375,0.015625,0.0234375,0.0234375,-0.015625,-0.0078125,0,0,-0.015625,-0.0234375,0.015625,0,-0.03125,0.0234375,-0.0234375,0,0.015625,0,-0.015625,0.0078125,0,0,-0.0078125,-0.0078125,-0.0078125,0,0.0078125,0.0078125,-0.0234375,0.015625,0,-0.03125,0.015625,-0.03125,0.03125,0,-0.0390625,-0.0078125,0.0234375,0,-0.0234375,0,-0.0078125,0.0390625,-0.0078125,-0.015625,0,-0.0234375,-0.015625,-0.0234375,-0.0234375,-0.046875,0,0.0234375,-0.03125,-0.0390625,0.046875,0.0078125,-0.0078125,-0.0234375,-0.03125,0.0078125,0,-0.0078125,-0.0078125,-0.0234375,0.0078125,0,0,-0.015625,-0.0234375,-0.015625,0.0234375,0.0234375,-0.0234375,0.03125,0.0390625,0.0078125,-0.0234375,0.046875,0.0078125,-0.0078125,0.03125,-0.0234375,-0.0390625,0.0078125,0.0078125,-0.03125,-0.046875,-0.0390625,0.046875,0.0078125,-0.0390625,0.0546875,0,-0.0234375,-0.0234375,-0.0078125,-0.0234375,-0.015625,0,-0.046875,-0.0078125,0.0546875,0.0078125,-0.0390625,0.0625,0.0546875,0,-0.0234375,0,0,0.0078125,0.0078125,-0.03125,-0.046875,-0.015625,0.0390625,0.0390625,0.0078125,0.0234375,0.0625,-0.0390625,-0.015625,-0.0234375,-0.03125,-0.03125,-0.046875,-0.015625,-0.0546875,-0.0390625,-0.0234375,-0.046875,-0.015625,0,-0.03125,-0.015625,-0.0078125,-0.015625,-0.03125,0.046875,0.0078125,0.03125,0.0234375,-0.03125,-0.0390625,-0.015625,0.015625,0.0078125,-0.015625,-0.0625,-0.0234375,0.015625,0.015625,-0.0078125,-0.015625,-0.0078125,0.046875,0.03125,0.0078125,-0.0390625,0.0078125,-0.0234375,-0.078125,-0.0078125,-0.0234375,0.03125,0,0.0234375,0,0,0.0234375,-0.0078125,-0.015625,0,-0.0078125,0,-0.03125,0.0390625,0.0390625,0.015625,-0.046875,-0.0078125,-0.0078125,-0.0078125,0.046875,-0.0390625,0.0390625,0.0078125,-0.03125,-0.015625,-0.015625,0.03125,0.015625,-0.0390625,0.0625,-0.0390625,-0.0234375,0.0078125,0.03125,-0.0546875,-0.046875,0,0.046875,0,-0.0078125,0,0,-0.0078125,0.015625,-0.0078125,0,0.015625,0,-0.0234375,0.015625,0.0546875,-0.015625,0.015625,0.0546875,-0.0546875,0,0.1015625,0.0390625,0.015625,-0.0546875,-0.0625,0.0390625,-0.0703125,-0.0078125,0,0.0078125,-0.0390625,-0.0546875,0.203125,-0.046875,0.0390625,-0.1328125,0,-0.0546875,-0.0234375,0.03125,-0.0078125,-0.0546875,-0.0546875,-0.03125,0.03125,0,-0.015625,0.0859375,-0.0703125,-0.0390625,-0.046875,-0.046875,-0.015625,-0.015625,-0.0234375,0.0390625,0,-0.03125,0.015625,0.046875,-0.0703125,0.0078125,-0.0546875,-0.0078125,0.03125,0.03125,-0.015625,0.0078125,0.0625,-0.03125,0.0078125,0.0234375,-0.0234375,-0.0234375,-0.0078125,-0.0703125,-0.0078125,0.0078125,0.046875,0.0078125,-0.0078125,0.0390625,0.0234375,0.0390625,-0.0546875,-0.0078125,-0.0546875,-0.015625,0.0078125,0.0234375,-0.0703125,0.0546875,0.0625,0.046875,-0.0078125,-0.0234375,-0.0859375,-0.0390625,-0.0234375,0,-0.0703125,-0.015625,0,-0.0078125,0,0.0078125,-0.0078125,-0.0078125,0.0078125,0.0078125,-0.0078125,-0.0078125,-0.015625,0.0078125,-0.0390625,-0.03125,0.0234375,0,-0.015625,-0.03125,0.0625,0.046875,-0.0859375,0.0703125,0.046875,-0.015625,-0.0390625,0.0390625,0.078125,-0.0390625,-0.03125,0.0390625,-0.0078125,0.03125,-0.0078125,-0.0390625,0.015625,0.0859375,-0.0546875,-0.0234375,-0.0390625,0.015625,0.03125,-0.0234375,-0.015625,-0.0390625,0.0078125,0.0546875,0.046875,-0.015625,-0.0546875,-0.109375,0.046875,0.078125,-0.015625,-0.0390625,0.0703125,0,0.046875,-0.0625,-0.015625,-0.0078125,-0.0625,0.015625,0,-0.0390625,-0.046875,0.046875,-0.0625,0.0859375,0,0.015625,0.0625,0.0703125,-0.015625,-0.0234375,0.03125,-0.0390625,-0.0078125,0.03125,0,0.015625,0.015625,-0.03125,0,0.03125,-0.0390625,-0.0390625,-0.015625,0.015625,0.0625,-0.0234375,0.0390625,0.046875,0.0078125,-0.015625,-0.03125,0.03125,0.0703125,0.0234375,-0.015625,-0.09375,-0.046875,0.0390625,0.1171875,0.015625,0.0078125,0.0234375,0.0546875,0.0078125,0.0234375,0,-0.015625,0.0625,0.03125,0.0625,-0.0859375,0.078125,-0.0546875,0.046875,-0.0390625,-0.03125,0.0625,-0.0625,0.03125,0.0703125,-0.046875,0.0234375,0.046875,0,0.015625,-0.046875,-0.03125,0.0078125,-0.0078125,0.015625,0,-0.0390625,-0.0390625,-0.046875,-0.0390625,-0.1015625,-0.0625,0.0546875,0.0546875,0.0625,0.015625,0,0.03125,0.03125,-0.0234375,-0.0234375,-0.046875,0.046875,-0.015625,0,0,0,-0.0078125,0.0078125,0,0.015625,0.0078125,-0.0234375,-0.0390625,0.0078125,-0.0234375,-0.0234375,-0.0546875,0.046875,-0.03125,-0.015625,0.0234375,-0.0078125,-0.0390625,-0.0234375,0.0078125,0.0390625,0,-0.046875,-0.0546875,-0.015625,-0.046875,0.0078125,-0.0078125,-0.0078125,0,-0.015625,0,-0.0078125,0,0.015625,0.0078125,0.0078125,0.0078125,-0.0078125,0,0.0078125,-0.0078125,-0.078125,0.0078125,0.0078125,0.0078125,0.0234375,-0.0234375,-0.03125,0.0234375,0,-0.015625,-0.03125,-0.0390625,-0.0234375,0.03125,0.0625,0.0078125,0.0703125,0.015625,0.0546875,-0.046875,-0.0546875,0.046875,0.0078125,-0.0546875,-0.015625,-0.0625,0.0390625,-0.0625,-0.0234375,-0.0390625,0.1015625,-0.015625,-0.0546875,-0.0078125,-0.015625,0.0078125,0.0078125,0,0,-0.0546875,-0.0234375,0.1015625,0.0078125,-0.0234375,-0.015625,-0.015625,0.0234375,0.0390625,-0.015625,0.015625,0.0390625,0.0078125,-0.0078125,-0.0234375,-0.015625,0,0.03125,-0.015625,-0.046875,0.0078125,0.0078125,-0.0390625,0.0390625,-0.0078125,0,-0.0078125,-0.015625,-0.015625,-0.0234375,0.03125,0.0234375,0.015625,0.0390625,0,-0.0234375,0.015625,0.015625,0,0,0,-0.015625,-0.03125,-0.1015625,-0.03125,0.0859375,0.015625,-0.0546875,-0.0234375,-0.0078125,-0.015625,-0.0078125,0.0078125,0.015625,0.0078125,-0.0078125,-0.0078125,0.015625,0.015625,0,-0.0390625,0.0234375,0.0234375,0.0078125,0.0546875,-0.0078125,0.03125,-0.015625,-0.03125,-0.0078125,0.0546875,0.0234375,-0.03125,-0.0078125,0.03125,0.015625,0,-0.03125,0.0859375,0.0390625,-0.03125,-0.0234375,-0.03125,-0.0546875,-0.015625,0.0234375,-0.0078125,-0.015625,0.015625,0.09375,-0.0234375,-0.078125,0.0078125,0.0390625,-0.0625,-0.0390625,-0.0546875,0.0234375,0.03125,0.0234375,-0.0625,-0.1171875,0.109375,-0.046875,-0.046875,0.0625,-0.0546875,-0.0234375,-0.015625,-0.0234375,-0.015625,0.0234375,-0.03125,-0.0078125,-0.0390625,-0.0546875,-0.0546875,-0.015625,0,0.078125,0.046875,0.0859375,0.0078125,0.0078125,-0.0390625,0.046875,-0.0234375,-0.0234375,0.0234375,0.0625,0.03125,-0.0625,0,0.0390625,0.03125,-0.0390625,0.0234375,0.09375,0.015625,0.078125,-0.015625,-0.0078125,0.0390625,0.046875,-0.0625,-0.046875,-0.046875,-0.0078125,-0.0859375,0.09375,0.0390625,-0.0703125,-0.0390625,0.0859375,0.0234375,-0.0078125,-0.125,-0.0703125,0.015625,0.0234375,0.03125,-0.09375,-0.078125,0.078125,-0.0234375,0,0.078125,-0.0078125,-0.03125,0.03125,-0.046875,-0.125,0.03125,0.125,-0.03125,0,0.0546875,0.015625,-0.078125,-0.078125,-0.0625,-0.078125,-0.0546875,0.015625,-0.0390625,-0.03125,0.0234375,0.0078125,0.0078125,-0.03125,-0.0078125,0.0859375,-0.0234375,-0.0625,0.046875,0.015625,0.140625,0.046875,-0.046875,-0.09375,0.0390625,0,-0.015625,-0.03125,0,-0.0078125,0,0.0234375,-0.015625,-0.0078125,-0.0078125,-0.0078125,0.0078125,0.109375,0.0703125,-0.0078125,-0.0078125,-0.0546875,0.0234375,0,0.015625,-0.0234375,0.0234375,-0.03125,0.015625,-0.0390625,-0.0234375,0.0078125,0.015625,0.0703125,0,0.0625,0.015625,0.0234375,-0.0078125,-0.0703125,0,-0.046875,-0.0390625,0,-0.015625,0.015625,-0.0078125,0.0078125,0,-0.015625,0,0.0078125,0.0078125,-0.0390625,0.0625,-0.09375,0.0234375,-0.0234375,0,0.046875,-0.0390625,-0.0078125,0.015625,-0.0078125,0,-0.046875,-0.140625,-0.0859375,-0.0078125,-0.015625,-0.046875,0.015625,0.0234375,0.0078125,0.0625,-0.03125,0.0078125,0,-0.0234375,-0.0078125,0.0234375,0.078125,0.046875,0.0390625,0.0390625,-0.0078125,-0.015625,-0.0234375,-0.0546875,-0.0390625,-0.0078125,-0.03125,-0.0390625,0.0078125,0.046875,-0.0625,-0.03125,-0.03125,0.015625,0,-0.0078125,0.03125,0.0078125,-0.03125,0.0234375,0.0078125,0.0078125,-0.0234375,0.015625,0.0078125,0.0078125,-0.0234375,0,0.0078125,0.0234375,0,0.015625,0.0390625,-0.0234375,0.0234375,0.046875,0.0078125,-0.03125,-0.015625,-0.0078125,0.03125,-0.078125,0.109375,0.09375,-0.0703125,0.0390625,-0.0078125,-0.0546875,-0.03125,0.1328125,-0.0546875,0,0.0234375,0.0078125,0.015625,0,-0.0234375,-0.015625,0.015625,-0.0078125,0.015625,-0.0078125,0.0234375,0.0234375,0,0,0.0078125,0,0.0078125,0.0078125,0.0078125,0,-0.0546875,0,0.015625,0.0078125,-0.046875,-0.0625,0.046875,0.1171875,-0.046875,0.0390625,0,-0.015625,-0.046875,0.0078125,-0.0625,-0.0390625,0.09375,-0.0234375,0,-0.046875,-0.03125,-0.0390625,-0.0390625,-0.078125,-0.0703125,0.140625,0.046875,0.109375,0.015625,-0.046875,0.03125,0.03125,-0.0234375,0.0390625,-0.015625,0.0078125,-0.03125,0.03125,0.03125,-0.0234375,0.0703125,0.0390625,0.0859375,-0.0234375,-0.0625,0.109375,-0.0078125,0.09375,0.03125,-0.1015625,0.1171875,-0.0234375,0.0234375,-0.0390625,-0.0390625,0,0.0546875,-0.0390625,0,0.0234375,-0.046875,-0.015625,0.03125,0.015625,-0.078125,-0.03125,0.0390625,-0.0234375,-0.0390625,0.0390625,-0.0234375,-0.0859375,-0.078125,0.03125,0.078125,0,0.015625,-0.03125,-0.0703125,0,0.0625,0.0234375,-0.0390625,-0.0234375,-0.0078125,0.1171875,-0.109375,-0.0234375,-0.0390625,-0.03125,0,-0.015625,-0.03125,-0.03125,0.046875,-0.0234375,0.015625,-0.03125,-0.0234375,-0.0078125,-0.015625,-0.0390625,-0.0546875,0.09375,-0.0234375,0.1015625,-0.0390625,-0.0625,0,0.0078125,0.0625,-0.0546875,0.078125,-0.046875,-0.0546875,-0.015625,-0.03125,0,0.015625,0.0234375,-0.03125,-0.0234375,0.0390625,0.0703125,-0.0390625,-0.046875,-0.1328125,0.015625,-0.0546875,-0.0546875,-0.046875,0.0078125,0.0078125,-0.078125,0.078125,-0.015625,0,-0.0703125,-0.078125,-0.0078125,0,0,-0.0078125,-0.015625,0,-0.015625,0.0390625,0,-0.03125,0.015625,-0.0390625,0,0,0.0078125,-0.078125,-0.0078125,-0.0390625,-0.0390625,0.0078125,-0.0390625,0.0078125,0.0078125,-0.0078125,0.03125,-0.0078125,0,0.015625,-0.0078125,-0.0390625,-0.078125,-0.0546875,0.0078125,0.0234375,0.015625,-0.0078125,-0.015625,0,0.0078125,0.0078125,-0.0078125,-0.015625,0.015625,-0.0078125,-0.0078125,-0.0390625,-0.03125,-0.0859375,-0.015625,-0.03125,0.046875,0.0390625,0.046875,0.03125,0.015625,-0.015625,0,0.046875,0.1484375,0,0,-0.0546875,0.0078125,-0.0078125,-0.0390625,-0.0234375,-0.03125,0.0234375,-0.0625,0.015625,-0.0625,0.0078125,0.0078125,0,-0.015625,-0.03125,0.0625,0.015625,-0.015625,-0.046875,0.0234375,-0.1171875,-0.0546875,-0.03125,-0.0234375,-0.0703125,0.0546875,0.1015625,0.0625,0.0546875,-0.03125,-0.03125,0.0234375,0,0,0,0.015625,0.0625,0.0234375,0.015625,0,-0.0234375,-0.015625,0.03125,0.03125,-0.03125,-0.015625,0.0078125,0.046875,-0.015625,0,-0.03125,-0.046875,0,0,-0.015625,-0.0390625,-0.0390625,-0.046875,0.0234375,-0.046875,-0.0703125,0.046875,0.0078125,0.0703125,-0.0625,-0.0078125,-0.03125,-0.0703125,0.0625,-0.015625,0.046875,0.015625,0.015625,-0.0078125,0.015625,-0.0078125,0.015625,-0.015625,0,-0.0078125,0.0078125,-0.0078125,-0.0234375,0.0234375,-0.0390625,-0.015625,-0.03125,-0.015625,-0.0078125,0.0234375,0,0.0390625,0.03125,0.03125,0,-0.0234375,0,-0.109375,-0.0078125,0,-0.046875,-0.0390625,0.015625,0,0,-0.03125,-0.0390625,-0.09375,0.015625,-0.0234375,0.046875,-0.109375,-0.03125,-0.0625,-0.0390625,0.0546875,-0.078125,0.109375,-0.0859375,0.015625,0,-0.0234375,-0.109375,0.0078125,-0.03125,-0.0234375,-0.09375,0.046875,0.0625,0.03125,0.0390625,-0.0546875,0.0234375,0.015625,-0.0546875,0.0234375,-0.0625,0.03125,0,-0.0390625,-0.03125,0.0078125,-0.0390625,-0.03125,0.0390625,-0.0703125,-0.0234375,-0.0234375,-0.0234375,-0.0546875,0,-0.046875,0.0546875,-0.015625,-0.0078125,0.0625,-0.0390625,0.1015625,0.0078125,-0.03125,0.03125,-0.0234375,0.0703125,-0.0703125,0.0390625,0.0703125,-0.0078125,-0.03125,0,0.0078125,-0.0390625,-0.046875,-0.015625,0.0078125,0.0859375,0.03125,0.0703125,0.03125,0.046875,-0.0546875,-0.1015625,-0.0390625,0.0234375,-0.078125,-0.046875,-0.0234375,-0.1171875,-0.0625,-0.015625,0.1015625,0.015625,0.0859375,-0.0546875,-0.015625,0.0078125,-0.1015625,0,0,0.03125,0.0625,0.0703125,-0.0078125,-0.015625,0.0390625,0.0625,0.015625,-0.0546875,0.0078125,-0.015625,0.046875,-0.078125,-0.0390625,-0.0078125,0.0234375,0,0.03125,0,-0.03125,-0.015625,-0.046875,-0.0234375,0,-0.0390625,0.0859375,0.0625,0.0703125,-0.0546875,-0.0078125,-0.015625,0.0078125,0.015625,0.0234375,-0.0078125,0.0078125,0.0078125,0,-0.015625,0.0078125,0.0625,-0.0078125,-0.109375,0.0625,0.015625,-0.0234375,0.0625,-0.0234375,-0.0078125,0.0234375,0.0390625,-0.03125,-0.0625,0,-0.015625,0.0546875,0.0390625,0.0390625,0.109375,-0.0078125,-0.015625,-0.0625,-0.0078125,0.015625,-0.0625,0.0078125,0.0078125,0,0,0.0078125,0.015625,0.0078125,0,0.0078125,0.0234375,-0.0234375,0.0078125,0.0859375,-0.046875,-0.078125,0.0859375,0.046875,-0.03125,0.0078125,0.0390625,-0.0390625,0.0703125,-0.015625,0.0703125,-0.078125,-0.0625,-0.0625,0.03125,-0.0234375,-0.0234375,0.0078125,-0.1484375,-0.0078125,0.0078125,0.09375,0.03125,0.0234375,-0.03125,-0.0078125,-0.0078125,-0.0703125,0,-0.046875,-0.0234375,0.0703125,0,-0.0078125,-0.0546875,-0.0078125,0,-0.015625,0,0.0546875,-0.0546875,-0.0234375,-0.046875,-0.046875,-0.0390625,0.109375,0.0234375,0.03125,0.0703125,0.0390625,-0.0234375,-0.0078125,0.015625,0.046875,-0.0390625,0.0234375,-0.0234375,-0.0234375,-0.015625,0.015625,0.046875,-0.03125,0.046875,-0.015625,-0.0234375,-0.0078125,0.015625,0.078125,0.015625,0.0390625,0.09375,-0.0234375,-0.046875,-0.0703125,-0.109375,0.09375,-0.0078125,0.015625,-0.0390625,0.0625,-0.0078125,0.0625,0.0859375,-0.015625,-0.0546875,0,-0.015625,-0.0078125,0,-0.015625,-0.0078125,-0.015625,0,0,-0.0078125,0,0.0234375,-0.0390625,-0.015625,0.03125,-0.015625,-0.03125,-0.0234375,-0.046875,-0.0078125,-0.0234375,-0.015625,-0.0390625,0.0234375,0.0703125,-0.046875,0.0078125,0.0390625,-0.0703125,0.015625,0.0078125,-0.0078125,-0.0234375,-0.0546875,0.0234375,0.078125,0.046875,0.1015625,0,0.015625,-0.0234375,-0.015625,-0.0234375,-0.0078125,0.0546875,0,-0.0234375,0.0078125,0.03125,-0.0390625,-0.015625,0.015625,-0.0078125,-0.0859375,-0.0390625,0,-0.03125,-0.03125,-0.0546875,-0.046875,-0.0390625,0.0234375,-0.015625,0.0859375,0,0.0234375,-0.0234375,-0.0234375,-0.015625,-0.015625,0.046875,-0.046875,0.046875,-0.03125,-0.046875,-0.0234375,-0.03125,0.0234375,0.03125,0,-0.0078125,-0.0390625,-0.03125,-0.046875,-0.015625,-0.0625,-0.09375,-0.0546875,-0.0625,0.078125,-0.0546875,-0.015625,-0.0234375,-0.0078125,0.0625,0,0.1015625,0.0390625,0.0859375,0.0078125,0.015625,-0.0859375,-0.03125,0.046875,-0.03125,-0.0390625,-0.0390625,0.046875,0.1015625,0.03125,0.0859375,0.0078125,-0.015625,0.0390625,-0.0703125,-0.0703125,-0.0859375,-0.0625,-0.0078125,-0.0078125,0.015625,0.03125,-0.0625,-0.0234375,0.015625,-0.0390625,0.046875,0.0234375,0.015625,-0.015625,0.0078125,0.0546875,-0.0625,-0.03125,-0.0703125,-0.046875,-0.03125,-0.0625,-0.0390625,0.046875,-0.078125,0.109375,0.046875,0,0,-0.015625,-0.0390625,0.0078125,0.0390625,-0.03125,-0.0234375,-0.0234375,-0.0078125,-0.0234375,0.0078125,-0.0078125,-0.0078125,0,-0.0078125,0.0078125,0.0078125,-0.0078125,0,-0.03125,0.015625,0.046875,0.0546875,0.078125,0.0078125,0.015625,-0.03125,-0.0078125,-0.046875,-0.015625,0.03125,0.0234375,0.015625,-0.0234375,0.0078125,-0.0234375,0.0390625,-0.078125,-0.015625,-0.0625,-0.0546875,0.0625,0.0625,0.0390625,-0.0390625,0,0.015625,0,0.0078125,0.0078125,0,0,0,-0.0078125,0,0.0078125,-0.0234375,-0.0078125,-0.0390625,0.03125,0.0546875,0.015625,-0.0546875,-0.03125,-0.0390625,0.03125,-0.0546875,0.09375,0.0234375,-0.0390625,-0.03125,-0.015625,-0.0078125,0.0390625,-0.015625,-0.0234375,-0.015625,0.078125,0.0546875,-0.0078125,-0.078125,-0.046875,0.015625,0,-0.0078125,0.015625,0.0546875,0.0234375,0.0078125,-0.015625,0.015625,0.0078125,0,0.0078125,-0.078125,-0.0234375,0.0234375,0.0078125,0,-0.03125,-0.0234375,-0.0078125,-0.0234375,0.0234375,-0.015625,-0.0625,0.015625,-0.015625,-0.0078125,-0.03125,-0.0078125,0.0078125,0.0625,0.0078125,0,-0.03125,-0.03125,0,0.0078125,0.0390625,0,0.0625,0,0.0234375,-0.0234375,-0.0078125,-0.015625,-0.03125,-0.0390625,0.015625,-0.0703125,-0.0703125,0.0390625,-0.0234375,0.0078125,-0.046875,0.0078125,-0.0234375,0.0078125,0,-0.0078125,0.0390625,-0.046875,-0.015625,0,0.0078125,-0.015625,0,-0.0078125,0,0.0078125,-0.015625,-0.0078125,-0.0078125,0,0.015625,0.046875,0.0390625,0.0390625,-0.0625,0,-0.0078125,-0.03125,0,-0.0078125,-0.03125,0.0234375,-0.0078125,-0.0390625,-0.015625,-0.0078125,-0.015625,-0.03125,-0.0625,-0.0625,0.0703125,0.0234375,0.03125,0.0078125,-0.015625,-0.0078125,0.046875,0.0703125,-0.0234375,-0.03125,0.078125,-0.0234375,0,-0.03125,-0.0390625,-0.03125,-0.0078125,0.0078125,0.1171875,0.109375,-0.03125,-0.0078125,-0.03125,-0.03125,0.0234375,0.015625,-0.0234375,0.0078125,0.0078125,-0.0546875,-0.0234375,0,-0.0234375,-0.0078125,-0.03125,-0.0078125,0.125,0.0390625,-0.0234375,0.0234375,-0.0703125,0,0.0703125,0.0703125,0.0390625,-0.0234375,0,-0.046875,0.015625,0.015625,-0.015625,0.0703125,-0.0234375,-0.046875,0.0234375,-0.03125,0,0,-0.015625,-0.015625,-0.0078125,0.0078125,-0.03125,0.03125,0.1015625,0.015625,-0.046875,-0.0234375,-0.0078125,-0.078125,-0.0390625,0.0234375,-0.03125,-0.0546875,0.015625,-0.0546875,0,0.015625,-0.0390625,-0.015625,-0.0546875,-0.0078125,0.03125,-0.0078125,-0.0390625,-0.0078125,0.015625,-0.0625,-0.0390625,0.0625,0,-0.0625,-0.0234375,-0.0078125,-0.015625,-0.0078125,0,-0.015625,0,0.0703125,-0.0703125,-0.015625,-0.0703125,-0.0078125,-0.0078125,-0.0390625,0.0234375,0.0078125,0.015625,0,0.0390625,0.0625,0.0234375,0.03125,-0.0234375,0,-0.0546875,-0.0390625,0.0390625,-0.0234375,-0.015625,0.0078125,-0.0234375,-0.0078125,0.0078125,-0.015625,0.015625,-0.0078125,-0.0078125,-0.0078125,-0.0078125,-0.0078125,-0.015625,0.0390625,-0.0859375,0.015625,0.03125,0.0078125,-0.0625,-0.0234375,0.078125,-0.0390625,-0.03125,-0.03125,0.0546875,0.0625,-0.015625,-0.03125,0.0078125,-0.0234375,-0.0234375,0,-0.0078125,0.0390625,0.015625,0.03125,0.03125,-0.0234375,-0.03125,-0.0078125,0.0234375,0.0078125,-0.0078125,0.0078125,-0.0078125,0,0.0078125,0,-0.046875,-0.03125,-0.140625,-0.0390625,-0.015625,0.0234375,0.0078125,0.0078125,0.0234375,-0.0390625,0.0234375,-0.0625,0,-0.109375,-0.0703125,-0.0234375,-0.0546875,-0.0078125,-0.03125,0.0078125,0.0078125,-0.015625,0.015625,0.03125,-0.015625,-0.0390625,-0.015625,0.015625,0.0078125,0.0078125,-0.0078125,-0.0234375,0.0234375,0.0078125,0,-0.015625,-0.015625,-0.046875,-0.0234375,-0.0703125,-0.03125,0.0390625,0.109375,0.0703125,0,0,-0.0234375,-0.0390625,-0.0078125,-0.015625,0,-0.0078125,0.03125,-0.0234375,0.0078125,0,0.015625,-0.03125,0.015625,-0.0078125,0,-0.03125,-0.0078125,-0.0078125,-0.0234375,0,-0.015625,0.1171875,0.046875,-0.0546875,-0.0703125,-0.0078125,-0.0234375,-0.0859375,-0.0078125,0.046875,-0.078125,-0.0546875,0.1171875,-0.0390625,-0.015625,-0.0546875,-0.0390625,0.03125,0,0.0859375,0.0078125,0.046875,0.0078125,-0.03125,0,0.0078125,-0.0078125,0.015625,0,-0.015625,-0.015625,0.015625,0.015625,0.0078125,0.015625,-0.0546875,-0.046875,-0.0234375,-0.0625,-0.0234375,-0.0234375,-0.03125,0.0234375,0.0078125,-0.0390625,0.015625,-0.0078125,0.0234375,0.0390625,-0.0078125,0.03125,-0.0546875,-0.0234375,-0.0234375,-0.078125,0.015625,-0.03125,-0.015625,-0.0078125,0.015625,-0.0234375,-0.015625,-0.0234375,0.046875,-0.015625,0.0625,-0.0546875,-0.0078125,0.0078125,-0.015625,-0.0078125,-0.0078125,-0.0078125,-0.0078125,0,0.0078125,0.0078125,-0.0234375,0.0078125,-0.0390625,0.015625,0.015625,0.0390625,0.015625,-0.0234375,0.0234375,0.0859375,0,-0.03125,0.0703125,-0.0625,0.0546875,-0.0703125,-0.03125,0.015625,0.0625,0,-0.015625,-0.0078125,-0.0078125,-0.0390625,-0.0390625,0.0234375,0.0703125,-0.015625,-0.0546875,-0.046875,0,0.0625,0.0078125,0.0625,0.0546875,-0.0390625,0.0078125,-0.0078125,0.046875,-0.046875,-0.0390625,0.078125,-0.0546875,-0.0625,-0.03125,-0.0078125,0.0546875,-0.0234375,0.0625,-0.0703125,-0.0390625,0.0390625,-0.0234375,-0.0703125,-0.03125,0.0078125,0.0234375,0,-0.078125,-0.0234375,0,0.046875,0.0078125,-0.0234375,-0.0546875,-0.0234375,-0.0234375,0,0.015625,0.0390625,0.0546875,0.0390625,0,0,0.03125,0,-0.03125,0.0625,-0.0234375,-0.03125,-0.015625,0.0234375,0.09375,0.0390625,0.0625,-0.015625,-0.015625,-0.0234375,0.0078125,-0.0859375,0,0.0078125,-0.0390625,-0.046875,-0.0390625,-0.0390625,0,0,-0.0078125,-0.03125,0,0.0078125,0,-0.0078125,-0.0078125,0.0078125,0.015625,0,0,-0.0546875,0,0.046875,-0.0234375,-0.03125,-0.015625,0.0390625,0.015625,-0.0703125,0.03125,0,0,0.046875,0,-0.0546875,0.0234375,0.0234375,-0.0546875,0.0234375,0.0234375,-0.0234375,-0.0390625,0.0078125,-0.0546875,0.0625,0.015625,0.0390625,-0.015625,0.0078125,0,-0.0078125,0,-0.015625,0.0078125,0,-0.0078125,-0.0234375,0.0078125,-0.03125,-0.046875,0.0625,-0.0078125,-0.0234375,0.0390625,-0.0234375,-0.015625,0.046875,-0.046875,-0.0234375,-0.03125,0,-0.0078125,-0.0078125,0.0234375,0.0546875,-0.046875,-0.03125,0.0234375,-0.0078125,-0.046875,0.03125,-0.109375,0,0.0078125,-0.0078125,-0.015625,-0.0078125,-0.0078125,-0.0078125,-0.046875,-0.0625,-0.0078125,0.046875,0.03125,0.0078125,0,-0.0234375,0.0546875,-0.046875,-0.0234375,0.0234375,0.0390625,0.0703125,-0.015625,-0.03125,0.015625,0,-0.0234375,-0.0078125,0.015625,-0.015625,0,-0.0234375,-0.0234375,0,0.0078125,0.0078125,0.03125,-0.0078125,-0.015625,-0.0078125,0.0078125,-0.015625,0.0234375,-0.0078125,0.0078125,-0.015625,0.0078125,-0.046875,-0.0859375,0.0234375,-0.03125,-0.0078125,0,-0.03125,0.015625,-0.0234375,-0.0625,-0.03125,-0.0546875,0.0234375,0.0234375,-0.0234375,-0.0078125,0,0.0546875,0,-0.0234375,0.0078125,0.0078125,-0.015625,-0.015625,-0.0234375,-0.015625,0.015625,0,0.0078125,0.0078125,0,0.03125,0,0.03125,0.0703125,0,0.0703125,0.046875,-0.03125,0,0.03125,-0.0625,-0.046875,0.0078125,-0.0390625,-0.0078125,0.0546875,0.015625,-0.015625,-0.046875,0.03125,-0.0078125,0.0078125,-0.0390625,-0.03125,0.0546875,0,-0.03125,0.046875,-0.0390625,-0.0078125,0.015625,0,0.0078125,0.109375,0.015625,0.0078125,0.0234375,-0.046875,-0.0078125,-0.046875,0.03125,0.03125,-0.0234375,-0.0234375,-0.015625,-0.0390625,-0.03125,0.0390625,0.015625,-0.0234375,-0.078125,0.1484375,-0.0078125,-0.0234375,-0.0234375,-0.0234375,0.015625,0.03125,0.03125,0.046875,-0.0390625,0.0234375,-0.03125,0.0078125,-0.0390625,0.03125,0.0234375,-0.0234375,-0.015625,0.046875,0.0625,-0.0859375,-0.0078125,-0.0859375,0.0390625,-0.0625,0.015625,0.015625,0,-0.0234375,-0.0078125,0.0546875,0.0390625,-0.0078125,0.0078125,0.0078125,-0.046875,-0.0078125,0.046875,-0.015625,-0.1171875,-0.0234375,-0.015625,-0.0703125,0.0390625,0.046875,0.03125,0.0390625,0.046875,0,-0.0234375,-0.0390625,-0.015625,0.0078125,-0.0234375,0.1015625,-0.0390625,0.015625,0,0.015625,-0.0234375,-0.0078125,-0.015625,-0.03125,0.078125,-0.0625,-0.03125,0.0078125,0.0078125,0.015625,-0.03125,-0.0234375,-0.0546875,0.0703125,-0.0390625,-0.0625,-0.0234375,-0.0546875,0.0546875,-0.0546875,-0.0078125,-0.03125,0.0078125,-0.03125,0.0078125,0.0234375,-0.0390625,-0.03125,-0.0234375,0,-0.0078125,0.0078125,0,-0.0078125,0.0078125,0.0078125,-0.0078125,0.0078125,0.0078125,-0.0234375,-0.0078125,-0.0078125,0.015625,0.046875,-0.0078125,-0.0234375,-0.03125,-0.0234375,-0.046875,0.0390625,0.0625,0,-0.0625,0.03125,-0.0078125,-0.0234375,-0.015625,0.0234375,-0.0234375,0.125,-0.015625,-0.1171875,-0.046875,0.0546875,0.015625,-0.015625,0,0.0078125,0,0.0078125,0,-0.0078125,0,-0.0078125,0,-0.046875,-0.0703125,-0.0078125,-0.078125,0.03125,0.03125,-0.0234375,0.015625,-0.0234375,-0.0625,0.0234375,-0.0234375,0.1015625,-0.1171875,-0.0546875,-0.0078125,-0.015625,0,-0.0234375,0.1484375,0.015625,0,-0.046875,-0.0234375,0.0234375,0.015625,-0.03125,-0.0078125,0.0078125,-0.0078125,0.046875,0.046875,0.0078125,-0.046875,-0.0390625,0,-0.0390625,0.046875,-0.0078125,-0.078125,-0.0234375,-0.0390625,-0.015625,0.0078125,-0.0234375,0.015625,0.0234375,0.0078125,0.0078125,0.0234375,0.0234375,0,0.0234375,-0.015625,0.03125,-0.015625,-0.0234375,0.0078125,0.0234375,-0.03125,-0.0078125,-0.0078125,0.015625,0.0390625,0,-0.015625,-0.0703125,0.015625,-0.0234375,0.015625,-0.0390625,-0.0078125,0.0390625,0,0.0546875,-0.0078125,-0.0078125,-0.03125,-0.0234375,-0.0078125,-0.0234375,-0.0546875,0,0.046875,-0.0234375,-0.0390625,-0.03125,-0.015625,-0.0390625,0,0.0078125,-0.015625,0.0078125,0.0078125,0,0.0078125,-0.015625,0.0078125,0,0,-0.015625,-0.0234375,0.0234375,0.046875,-0.015625,-0.0078125,0,0.0078125,0.0625,-0.015625,-0.015625,0.0546875,0.03125,-0.0234375,-0.046875,0.0234375,-0.0078125,-0.0390625,-0.0390625,-0.0078125,-0.0234375,0,0.09375,-0.0234375,0.0078125,0,0.015625,0.015625,0.0078125,0.0234375,-0.0390625,-0.046875,-0.03125,0,-0.0078125,0.0234375,-0.03125,0.0859375,0.0625,0.0234375,-0.0234375,-0.0703125,-0.0625,-0.0078125,0.0234375,0.015625,-0.0703125,0,0.0859375,0.015625,0.0234375,0.015625,0.0078125,0,-0.0703125,-0.0703125,0.015625,0.03125,0.09375,0.046875,0.0078125,-0.0234375,-0.0390625,0.078125,-0.0703125,-0.0078125,-0.0625,0.0078125,-0.015625,0.0078125,-0.015625,0.03125,0.03125,0.0390625,-0.0078125,-0.03125,-0.015625,0.0234375,-0.0546875,-0.015625,-0.0078125,-0.0234375,-0.015625,0.0234375,0.015625,-0.0859375,-0.015625,-0.046875,0,0.0703125,-0.0390625,-0.0390625,-0.0546875,0.0234375,-0.078125,0.046875,-0.03125,-0.0546875,-0.0078125,0.015625,-0.0234375,-0.0078125,-0.03125,-0.0390625,-0.015625,-0.03125,-0.015625,0.0078125,0,0.0234375,-0.0546875,0.03125,0.0390625,0,-0.03125,-0.0234375,-0.0234375,-0.0078125,-0.046875,0.0390625,-0.0234375,0.03125,0.0078125,-0.0234375,0.015625,0.015625,0.03125,-0.0234375,0.03125,0.0546875,0.015625,-0.046875,-0.03125,-0.0234375,-0.0234375,0.0078125,-0.0234375,-0.0625,0,-0.0234375,-0.0078125,-0.0234375,-0.0546875,0,0,0,-0.0078125,-0.0078125,0,0,0,-0.015625,-0.0234375,0.1015625,0.03125,0.0703125,0.046875,-0.0390625,0.015625,-0.015625,-0.03125,0.0078125,-0.03125,-0.0078125,0.0390625,0.0703125,-0.015625,-0.015625,-0.015625,-0.046875,0.0390625,0.1015625,0.03125,-0.0078125,-0.0390625,-0.0234375,-0.078125,0.0234375,0,-0.0078125,-0.0078125,0,-0.0078125,0,0,0.0078125,0.0078125,0.0078125,-0.0390625,0.0546875,-0.03125,0.046875,0.0234375,-0.0390625,0.0078125,0.1015625,0,-0.015625,0.03125,0.015625,-0.0859375,0,-0.0234375,-0.03125,0.0078125,-0.015625,-0.0078125,0.0546875,-0.0078125,-0.0625,0.015625,-0.0078125,0.03125,0.015625,-0.015625,-0.046875,0,0,0,0.0390625,0.015625,-0.046875,-0.0390625,-0.0078125,-0.03125,-0.0234375,-0.0390625,0.0390625,-0.0078125,-0.03125,-0.0390625,-0.0390625,-0.03125,-0.0546875,-0.015625,-0.046875,-0.03125,-0.03125,-0.015625,0,0.0703125,0,0.0078125,0.046875,-0.015625,-0.0078125,-0.0078125,0,-0.0234375,-0.0546875,0.0234375,-0.0078125,0.015625,-0.0234375,-0.015625,0.0078125,0.015625,0,0.0234375,0.03125,-0.0390625,-0.0546875,-0.0078125,0,0.015625,0.0078125,0.078125,-0.03125,-0.03125,0.015625,-0.0078125,0,-0.0625,0.046875,0,0.015625,0.046875,0.0078125,0.0078125,-0.0078125,0.0078125,0,0,-0.0078125,0,0,0,-0.0234375,0,-0.0078125,0,0.0234375,0,0.015625,0.078125,0.0078125,0.0078125,-0.015625,0.015625,-0.0234375,-0.015625,-0.0234375,-0.0703125,-0.046875,-0.0234375,-0.0078125,-0.0234375,-0.015625,0.0234375,-0.0234375,-0.03125,0.046875,-0.015625,-0.015625,-0.0390625,-0.078125,-0.015625,0.03125,-0.0703125,-0.0078125,-0.0078125,-0.0390625,0,0.0546875,0.03125,-0.03125,-0.0078125,-0.015625,-0.0078125,0.0078125,-0.0234375,0.0234375,-0.0078125,-0.03125,0.0234375,0.03125,-0.0078125,-0.0546875,0.03125,0.046875,0,-0.0390625,-0.03125,-0.0078125,0.03125,-0.0390625,-0.0078125,0.109375,-0.015625,-0.03125,0.0234375,-0.0234375,-0.0078125,0,-0.015625,-0.015625,-0.015625,0.046875,0,-0.0390625,-0.03125,-0.0078125,0.0234375,0.0390625,-0.015625,-0.0703125,0.0078125,0.046875,0.0078125,0.015625,0.03125,-0.046875,-0.0390625,-0.03125,-0.0703125,0.015625,0.0390625,-0.0390625,0.046875,-0.015625,0.0390625,-0.015625,0.0078125,-0.015625,-0.015625,0.0625,-0.0234375,-0.0390625,-0.03125,0.0625,-0.0625,-0.0390625,-0.03125,-0.0390625,-0.03125,-0.0234375,-0.0078125,-0.015625,0,0.0859375,-0.0234375,-0.015625,0,-0.0234375,0.015625,0.0234375,0.015625,-0.0703125,0.015625,-0.0390625,0,-0.0078125,0.0234375,0,-0.0703125,-0.015625,-0.0625,0.0078125,-0.03125,-0.03125,0.03125,-0.015625,-0.03125,-0.046875,-0.0703125,-0.0078125,-0.0234375,-0.046875,-0.0078125,0.046875,0.09375,0.0078125,0.0078125,0.0078125,-0.0078125,-0.0078125,-0.0078125,-0.0078125,0.0078125,0.015625,-0.0546875,0.046875,0.0546875,-0.03125,0.0234375,-0.046875,-0.046875,0.015625,0.0234375,-0.0078125,0.0390625,0.078125,0.0390625,0.0546875,-0.0234375,-0.0390625,-0.015625,0.0859375,-0.0546875,0,-0.0390625,0.03125,0.046875,-0.0546875,0.0078125,0.0625,-0.0078125,0,-0.0078125,0.0078125,0,0.0078125,0,-0.0078125,-0.015625,-0.0078125,0.0078125,-0.0859375,0.078125,-0.015625,-0.015625,-0.0625,-0.0234375,-0.046875,0.0390625,0.03125,-0.046875,-0.015625,-0.015625,-0.046875,-0.0859375,0,0.03125,-0.0234375,-0.0078125,-0.015625,0,0.0703125,0.0859375,-0.0390625,-0.0078125,-0.0078125,-0.046875,0,0.0390625,-0.046875,-0.0390625,0.0390625,0.015625,0.0234375,0.0234375,-0.03125,0,0.0703125,0.0078125,-0.1015625,0.0078125,0.03125,0,0.0546875,0.0390625,0,0.0078125,-0.0078125,0.0078125,0.0078125,-0.03125,-0.0234375,-0.0546875,-0.0390625,0,-0.0234375,0.0390625,0.0390625,-0.0078125,-0.015625,-0.015625,0.0078125,0,0,-0.0234375,0,0,-0.015625,0.1640625,0,-0.03125,0.0078125,0.0234375,-0.0078125,-0.125,-0.0703125,0.0859375,0.078125,-0.046875,-0.09375,-0.0703125,-0.0078125,0.0234375,0.0234375,-0.03125,0.0234375,-0.0390625,-0.046875,-0.0078125,-0.046875,-0.0078125,-0.0234375,0.0078125,0.0078125,-0.03125,0.015625,-0.0078125,0.0078125,-0.0078125,-0.03125,0.015625,-0.0625,-0.015625,0.015625,-0.0234375,0.0390625,-0.0078125,0.015625,0.046875,0.0390625,0,-0.0078125,0.0078125,0,0,0,0.0234375,-0.0390625,-0.0546875,-0.03125,-0.015625,0.0078125,0.0078125,-0.0390625,-0.03125,0.015625,0.0390625,-0.015625,-0.015625,0.03125,0,0.0703125,0.015625,0.015625,-0.0078125,-0.03125,-0.0390625,-0.0390625,-0.03125,0.0234375,0,-0.046875,0.015625,0.03125,0.0078125,0.0390625,-0.09375,0.0234375,0,-0.046875,-0.0546875,0.015625,-0.0078125,-0.015625,-0.0390625,0.1640625,-0.0625,-0.046875,-0.09375,0.0078125,0.046875,0.0078125,-0.046875,-0.015625,0,0,0.0390625,0,-0.0390625,0.0859375,-0.0546875,-0.0390625,0.0078125,-0.0625,-0.0546875,0.0625,0.015625,0.03125,0.03125,-0.0390625,-0.0234375,-0.03125,-0.0234375,0.0859375,-0.1171875,0.0234375,-0.046875,-0.0390625,0.046875,0,0.0625,-0.09375,0.03125,-0.015625,0.0859375,0.078125,-0.09375,-0.0625,-0.0078125,-0.0390625,-0.0234375,-0.046875,0.0390625,0.0546875,0.078125,-0.0390625,0,-0.0625,0,0.09375,-0.078125,0,-0.109375,0.1015625,-0.0625,0.0703125,0.0546875,-0.0078125,-0.0234375,0.0078125,-0.0078125,-0.0390625,0,0.0546875,0.0390625,-0.0703125,-0.0234375,0.046875,-0.0625,-0.0390625,-0.046875,-0.0078125,-0.0625,0.078125,0.015625,0.0703125,-0.0234375,0.0078125,-0.0078125,-0.0078125,-0.0390625,-0.046875,-0.0234375,-0.015625,0,-0.015625,0,0.015625,0,0.0078125,0.0078125,0,-0.0390625,-0.0234375,-0.0625,-0.0078125,-0.078125,-0.0703125,0.03125,0,0.015625,0,-0.03125,-0.0390625,0.0078125,0.0078125,-0.0234375,-0.03125,0,0.0078125,0.0078125,0.0234375,-0.046875,-0.078125,0.0078125,-0.015625,-0.03125,0.015625,-0.0078125,0.0078125,0.015625,0.0078125,0,-0.0078125,0,-0.0078125,0.0078125,-0.0078125,-0.0625,-0.0546875,-0.0703125,-0.015625,0.015625,-0.0625,-0.0234375,-0.0078125,0.015625,0.0078125,-0.015625,0,-0.015625,0.0390625,0.0703125,-0.0078125,0.0234375,0.0234375,-0.03125,0,0.0078125,0.0390625,0.0390625,0.0703125,0.0390625,-0.0234375,0.0078125,-0.03125,0.0078125,0.0234375,-0.0078125,-0.03125,0.0390625,0,0.0234375,0.0234375,0.0390625,-0.0546875,-0.015625,0,0.046875,0.015625,-0.0234375,-0.015625,-0.0078125,-0.0078125,0.03125,-0.0234375,-0.0234375,0.0078125,-0.0234375,-0.015625,-0.015625,0,-0.015625,-0.015625,0.0390625,-0.0078125,-0.0390625,0.0078125,-0.0234375,-0.0078125,0.0234375,0,0,-0.0078125,-0.03125,-0.046875,-0.0078125,-0.0234375,0.015625,-0.015625,0.03125,-0.0546875,0.03125,0.0234375,-0.0078125,0.0703125,-0.0234375,-0.0234375,-0.0546875,0.046875,-0.0234375,-0.0390625,-0.0234375,0.0234375,-0.03125,-0.03125,0.0078125,0,-0.0078125,-0.0078125,0.0078125,0.0234375,0,-0.0078125,-0.015625,0.0078125,-0.015625,-0.015625,0.03125,0.0390625,-0.015625,-0.015625,-0.03125,-0.0234375,-0.0078125,0.015625,-0.0390625,0.03125,0.03125,-0.0234375,0.015625,-0.0078125,0.0546875,0,0.0078125,-0.03125,0.0390625,0,-0.03125,0.015625,0,-0.0078125,-0.0546875,-0.0078125,-0.0078125,0.09375,-0.03125,0.015625,0.0703125,-0.0859375,-0.046875,-0.0390625,-0.03125,-0.015625,-0.0234375,0,0,-0.0078125,0,0,0.0390625,0.0078125,-0.0859375,0.109375,-0.0625,-0.0078125,0.0078125,-0.0546875,0.0625,-0.0234375,-0.0078125,0.125,-0.015625,0.046875,-0.0546875,-0.015625,-0.078125,-0.0546875,-0.015625,0,-0.015625,0.015625,0.0078125,-0.046875,0,-0.0390625,-0.0078125,0.0390625,0.015625,0,0,-0.0546875,0.0390625,0.0078125,0.0390625,0.046875,0.0625,0.0703125,-0.03125,-0.015625,0.03125,0.015625,0.0234375,0.0234375,-0.0625,-0.0546875,-0.046875,0.0625,-0.0234375,0.0390625,0.0078125,0.0234375,0.0234375,-0.046875,0.03125,-0.0234375,0.03125,0,0.0078125,-0.0234375,-0.0546875,-0.015625,0.0078125,0.0234375,0.0078125,0.0078125,-0.0234375,-0.0078125,0,-0.0546875,0,0.046875,-0.046875,0.0546875,-0.046875,0.140625,-0.03125,-0.0390625,-0.0390625,-0.0390625,0.0078125,-0.03125,-0.0390625,0.1015625,0.0390625,-0.0234375,-0.046875,-0.046875,0.0546875,0.0078125,0.0234375,-0.0546875,-0.03125,-0.0546875,-0.0078125,-0.0625,0,-0.0078125,-0.046875,0.1015625,0.0234375,0.0078125,0,0.0078125,0,0.0078125,0.0078125,-0.015625,0,-0.0078125,-0.0546875,0.046875,0.046875,-0.0625,-0.0234375,0.0390625,-0.0234375,0,-0.0234375,0.0078125,0.0625,0.0078125,-0.0390625,-0.03125,-0.03125,-0.0234375,-0.0234375,0.0078125,0.1015625,0.0546875,-0.046875,-0.0078125,-0.0546875,-0.0234375,0.0078125,-0.0078125,0.03125,0,-0.0078125,0,0,-0.015625,0.0078125,-0.0078125,-0.0078125,0.0078125,0,0.046875,0.0078125,0,0.0390625,-0.046875,-0.015625,-0.03125,0.0234375,0.0390625,-0.046875,0.0546875,-0.0546875,-0.0703125,-0.0390625,-0.03125,-0.0234375,-0.0390625,0.171875,0.015625,-0.046875,-0.03125,0.015625,-0.0390625,-0.015625,-0.03125,-0.0078125,-0.0078125,0.0078125,-0.015625,-0.03125,0.0234375,0.0234375,-0.046875,-0.015625,-0.0078125,-0.0703125,0.0546875,0.015625,0.0625,0.015625,-0.0390625,-0.0546875,-0.0234375,-0.03125,0.0625,0,-0.0546875,0,0.0390625,-0.0078125,0.015625,0.0078125,0,0.03125,-0.015625,-0.015625,-0.0078125,-0.015625,0.0078125,-0.015625,-0.015625,-0.0390625,0,0.0234375,-0.0078125,-0.046875,-0.0078125,0.015625,0.03125,-0.015625,-0.0234375,0,-0.046875,0,0.015625,-0.03125,-0.046875,-0.0390625,0.0546875,-0.015625,0.046875,0.046875,-0.0625,-0.0859375,-0.046875,0,0.0390625,-0.015625,0,0,-0.0078125,-0.0078125,0.0234375,0,0.0078125,-0.0078125,-0.0078125,0.0234375,0.0078125,0.0078125,0.0078125,-0.0390625,0.0390625,-0.03125,-0.0234375,0.0078125,0,-0.0390625,0.015625,0.0625,-0.0390625,0.0234375,0.0078125,0,-0.0078125,-0.015625,0.0625,0,-0.0234375,0.015625,-0.046875,-0.0234375,-0.0078125,0.015625,0.015625,-0.046875,0.046875,0.0625,0.046875,-0.0234375,-0.0546875,-0.015625,-0.0234375,0,0.0078125,-0.0390625,0,-0.1015625,0.0078125,0.0078125,-0.015625,0.015625,0.0234375,-0.0234375,0.0234375,-0.0546875,0.0546875,-0.0859375,-0.0234375,0.015625,0.0078125,0.03125,0.171875,-0.0390625,0.0078125,-0.0078125,-0.0703125,-0.03125,-0.0078125,0.015625,0.015625,0,0.0234375,-0.0390625,0.0859375,0.0078125,-0.0625,-0.0859375,-0.015625,-0.03125,0,-0.0859375,0,0.09375,-0.140625,0.0234375,0.0234375,0.0078125,-0.015625,-0.0078125,0.0078125,0.0625,-0.03125,0,-0.0078125,-0.0234375,0.0078125,0.046875,-0.0078125,0.046875,-0.046875,-0.0234375,-0.015625,0.0546875,0.03125,0,-0.0234375,0.0234375,-0.0234375,0.0859375,0.0703125,-0.046875,0.046875,-0.015625,-0.046875,-0.015625,0.046875,0.0625,0.03125,0.046875,0.0078125,-0.015625,-0.046875,-0.03125,-0.046875,-0.0078125,-0.015625,-0.0078125,0.0390625,-0.0234375,0.015625,-0.03125,-0.046875,0.0078125,-0.0546875,-0.0390625,0.0078125,-0.0078125,-0.03125,-0.0234375,0.0078125,0.0078125,0.03125,-0.046875,0.0234375,-0.0234375,-0.046875,-0.0078125,-0.03125,0.0625,0.046875,0,-0.0078125,-0.015625,0.0078125,-0.0078125,-0.0078125,-0.0078125,0,0.0078125,-0.0078125,0.0234375,-0.046875,-0.0625,-0.0234375,-0.0625,0.0625,0.125,0.015625,-0.046875,-0.0390625,0.0625,-0.0703125,0.0546875,-0.0546875,-0.0390625,0.0234375,0.0625,-0.015625,0.0546875,-0.03125,-0.0546875,-0.0703125,-0.03125,-0.0625,-0.0390625,-0.09375,-0.0703125,0,0.0078125,0,0,0,-0.0078125,0.0078125,0,0,-0.1171875,0.0234375,-0.0546875,-0.0078125,0.0390625,-0.09375,-0.0078125,0.078125,-0.046875,-0.0390625,-0.046875,0.0390625,0.03125,-0.0625,-0.0234375,-0.03125,0.015625,-0.0078125,0.0390625,0,-0.015625,-0.0390625,-0.078125,-0.015625,-0.0078125,-0.03125,-0.1015625,-0.0390625,-0.0390625,0.015625,0.046875,0.015625,0.0390625,0,0,-0.0078125,-0.0625,0.0078125,0.015625,-0.0078125,0.0546875,-0.03125,-0.0078125,-0.015625,0.015625,-0.015625,-0.0234375,0.015625,-0.0234375,-0.015625,0,-0.0234375,-0.0390625,0.0078125,-0.015625,-0.0078125,0.0078125,0.0546875,-0.0234375,-0.015625,-0.0234375,-0.03125,0.0078125,0.0078125,0.0234375,0,0.0078125,-0.0234375,0.0625,-0.03125,0.0390625,-0.0078125,-0.046875,-0.0390625,0,0.078125,0.0859375,-0.03125,0.0078125,-0.0390625,0.0390625,-0.0625,0.0078125,0,-0.0234375,-0.0078125,-0.03125,0.03125,-0.0703125,0.03125,0,0,0.0234375,0.015625,0.0390625,0.0078125,0,0.015625,0,0,-0.0078125,-0.0390625,0.015625,0.0078125,-0.046875,0.0390625,0,-0.0703125,-0.015625,0.0390625,-0.09375,-0.015625,0.046875,-0.109375,-0.078125,0.109375,-0.0234375,0.015625,-0.03125,0.015625,0,-0.0234375,-0.03125,-0.0234375,-0.015625,-0.0078125,0.03125,0.0546875,0.015625,0,0,0.0234375,-0.0390625,-0.0625,0.0390625,-0.125,-0.0703125,-0.0078125,0.0234375,-0.046875,-0.0546875,0.15625,0,-0.0625,-0.015625,-0.078125,-0.03125,-0.0625,-0.0390625,0.0625,0.0078125,0.0234375,0.015625,0,-0.03125,0.078125,-0.046875,-0.0390625,0.0859375,0.09375,0.1328125,0.0078125,-0.0234375,-0.0546875,-0.03125,-0.0234375,-0.0234375,0.015625,0.078125,-0.0234375,-0.015625,-0.0234375,-0.078125,-0.03125,-0.03125,0.0703125,0.0234375,0.015625,0.046875,0.046875,0.015625,0.0546875,0.0390625,-0.0234375,-0.0625,0.0078125,-0.0390625,0.0234375,0.0078125,0.109375,-0.0234375,0.0234375,0.0078125,-0.015625,0.0703125,-0.03125,-0.03125,0.0234375,0.046875,0,0.0078125,-0.046875,0.09375,0.0703125,-0.09375,0.0703125,0.0234375,-0.0078125,-0.0234375,0.0625,0.0703125,0.03125,0.0546875,-0.0078125,0.03125,0.015625,0.0625,0.015625,-0.015625,-0.046875,-0.1015625,0.0390625,0.03125,0,0.0546875,0.0078125,-0.03125,0.0234375,-0.03125,-0.03125,-0.078125,0,-0.0859375,0.0078125,0.03125,0.03125,0.0078125,-0.0390625,-0.0078125,-0.0078125,0,-0.0390625,-0.015625,-0.0078125,-0.0078125,0.0078125,0.0078125,0.0234375,0.0078125,0.0078125,0,-0.0078125,-0.03125,-0.0390625,-0.015625,-0.015625,0.015625,0.0078125,0.03125,-0.0078125,0.0078125,-0.03125,-0.015625,-0.015625,0.0078125,0,-0.0234375,-0.015625,-0.0390625,-0.015625,-0.0390625,-0.015625,0.0078125,0.03125,-0.0234375,-0.015625,-0.0234375,0.03125,0,0,0.0078125,0.0078125,0.0078125,0.0078125,-0.0078125,0.0078125,-0.0078125,0,0,0.0234375,-0.0234375,-0.0078125,0.0703125,-0.015625,-0.015625,0.0390625,0.0078125,-0.015625,-0.0546875,0.0078125,0,-0.0078125,0.0078125,-0.015625,0.015625,0,0.015625,-0.0625,-0.015625,0.0546875,0.03125,-0.03125,-0.03125,-0.0234375,-0.015625,-0.03125,0.0078125,0.0078125,0.03125,-0.0078125,0,0,-0.0234375,0.015625,-0.0234375,-0.015625,-0.015625,-0.0390625,0,-0.015625,-0.015625,0,-0.0234375,-0.0078125,-0.03125,-0.0078125,0.0078125,-0.015625,-0.0234375,-0.0078125,-0.015625,0.0078125,0.0078125,0,-0.015625,0.0234375,0.0546875,0,-0.015625,0.015625,-0.0078125,0.03125,0.015625,-0.0078125,0.046875,0,0.0078125,-0.0078125,0.0234375,0.0078125,-0.03125,0.03125,0,-0.015625,-0.03125,0,-0.0390625,-0.03125,-0.015625,0.03125,0.0625,-0.0078125,0,-0.03125,-0.0234375,-0.015625,-0.015625,-0.0078125,0,-0.0078125,-0.0078125,0.0078125,0.0078125,-0.015625,-0.015625,0.0078125,0.0078125,-0.03125,-0.0546875,0.0078125,0.03125,0.046875,0.0078125,0.015625,-0.015625,0.0078125,-0.0703125,0.0078125,-0.0234375,-0.015625,0.03125,-0.0078125,-0.0078125,-0.015625,0,0.03125,0,-0.0234375,0,-0.0390625,0.015625,-0.0390625,0.03125,-0.0078125,-0.0078125,-0.0078125,0,0.0234375,0,0.015625,0,0.0078125,-0.0078125,-0.046875,0.0078125,-0.0234375,0.0703125,-0.0234375,-0.0390625,-0.0234375,0.0078125,-0.0078125,0.03125,-0.0078125,-0.0078125,-0.0390625,0.0078125,0,-0.0078125,-0.0234375,-0.03125,0.0390625,-0.03125,-0.03125,0.0078125,0.0859375,0.0078125,-0.0234375,0,-0.046875,-0.0859375,-0.03125,0,0.0234375,0.0390625,-0.0078125,0.0390625,-0.0078125,-0.0078125,-0.0234375,-0.015625,-0.0078125,-0.046875,-0.015625,-0.015625,-0.0234375,-0.0078125,-0.0234375,0.0234375,0.015625,0,0.0078125,-0.0390625,0,-0.015625,-0.0234375,-0.0078125,0.046875,0.046875,0,0.046875,-0.015625,0.015625,-0.0390625,-0.0546875,-0.0234375,-0.03125,-0.015625,-0.015625,0,0,0.0390625,-0.0234375,0.03125,0,-0.03125,-0.0078125,-0.015625,-0.046875,0.046875,0,-0.0390625,-0.0546875,0.0078125,-0.03125,-0.015625,-0.0078125,-0.0078125,0,-0.0078125,-0.015625,0.0234375,0.0234375,-0.0546875,-0.0234375,-0.015625,0.015625,0,0,-0.0234375,-0.03125,0.015625,-0.0078125,0.0703125,0.1328125,-0.0546875,0.015625,-0.03125,-0.0078125,0.0703125,0.0234375,-0.0078125,0.0078125,0.0078125,0,-0.0078125,0,-0.015625,0,-0.0078125,-0.0078125,-0.0703125,-0.046875,-0.0390625,0.046875,0,0.03125,0.0546875,-0.0234375,-0.0234375,-0.015625,0.015625,-0.0078125,-0.015625,-0.0234375,-0.015625,0.0703125,0.046875,0.0078125,-0.0390625,-0.0546875,-0.0234375,0.0234375,-0.046875,0,0.0078125,0.03125,0.015625,0.0078125,0.015625,0,-0.0078125,0,-0.0078125,0.0078125,0,-0.0234375,-0.0546875,-0.0078125,0,-0.0390625,-0.046875,-0.0234375,0.015625,0.03125,0,-0.0390625,0.125,-0.015625,-0.1015625,-0.015625,0,-0.015625,0.0234375,-0.0078125,-0.0234375,-0.046875,-0.0234375,0.03125,0.0390625,-0.0546875,0.0078125,-0.046875,-0.0078125,-0.0390625,0.015625,-0.0625,0.0625,0.0390625,0.015625,-0.015625,-0.015625,-0.015625,-0.03125,0,0.0390625,-0.015625,-0.03125,-0.0390625,0.0625,-0.0078125,-0.0078125,0.015625,-0.015625,0,-0.03125,-0.0234375,-0.0234375,-0.0546875,-0.0234375,-0.0078125,-0.03125,0,0,0.015625,0,0.0078125,0,0,0.0078125,0.0078125,0.0078125,0.0078125,-0.0078125,-0.0234375,0,0.0390625,0.09375,-0.0234375,-0.0078125,0.0390625,-0.0390625,0.015625,-0.0625,-0.015625,-0.0546875,0.140625,0,-0.078125,-0.0546875,-0.0703125,-0.0625,0.0234375,0.0234375,0.0625,-0.0078125,0,-0.015625,-0.015625,0,-0.0078125,-0.015625,0.0078125,-0.0078125,0.015625,0,0.0078125,0.0234375,0.0078125,-0.015625,-0.03125,-0.0390625,0.0078125,-0.0234375,-0.015625,-0.046875,-0.0859375,-0.046875,0.0390625,-0.03125,-0.0234375,-0.015625,-0.015625,-0.015625,0.015625,-0.0234375,-0.0078125,-0.015625,-0.0703125,0.015625,-0.0703125,0.0859375,0.015625,0.03125,-0.1171875,-0.0546875,0,-0.046875,-0.0078125,0.0234375,0.1796875,-0.0078125,0,0.0390625,-0.0546875,0.0390625,-0.0546875,-0.03125,0.0078125,-0.046875,-0.0078125,0.03125,-0.0625,-0.0234375,0,-0.0859375,-0.0078125,-0.0078125,-0.0234375,-0.0078125,-0.0625,0.015625,-0.015625,-0.03125,0.046875,0.0078125,-0.0390625,-0.1484375,-0.0078125,0.0234375,-0.0078125,-0.0546875,0.0078125,-0.0625,-0.0625,-0.03125,0.0078125,-0.0078125,0.03125,-0.0390625,0,-0.0625,-0.0703125,-0.0078125,-0.03125,0,0.015625,-0.046875,0.03125,0.015625,-0.015625,-0.0234375,0,0.0234375,0.0234375,-0.0234375,-0.1171875,-0.0625,-0.0234375,0.1328125,0.046875,0.015625,0.0625,0.0078125,-0.015625,-0.0625,-0.0390625,0,-0.046875,0.015625,0.015625,-0.0546875,-0.0234375,-0.0078125,-0.0234375,-0.078125,0.0390625,-0.03125,-0.0078125,0.0234375,-0.0390625,-0.109375,-0.0078125,-0.015625,-0.046875,0.046875,-0.0078125,-0.03125,0.0078125,0.015625,0.0625,-0.0234375,0.03125,0.09375,-0.0078125,0,0.0703125,0.0078125,-0.015625,-0.0859375,0.03125,0.0078125,-0.0390625,-0.0078125,-0.0234375,-0.0234375,0.03125,-0.046875,-0.0234375,-0.015625,-0.0078125,0.0234375,0,0.015625,0.015625,-0.0078125,-0.0078125,-0.0078125,-0.1015625,-0.015625,-0.0625,0.015625,-0.0390625,-0.0390625,0.03125,0.015625,0,-0.0625,-0.0078125,-0.03125,-0.0078125,0.0859375,-0.0703125,0.03125,0.0078125,0.0234375,-0.0234375,-0.0703125,-0.046875,0.078125,-0.015625,0,-0.0625,-0.0546875,0,0.015625,0.0078125,-0.0078125,0.015625,0.0078125,-0.0078125,-0.0078125,0.0078125,0.0078125,-0.09375,0.1171875,-0.015625,0.0078125,-0.078125,-0.0390625,0.046875,-0.0078125,-0.015625,-0.0078125,-0.0078125,-0.0234375,-0.0078125,0.03125,-0.0078125,-0.046875,-0.0234375,0,0.0625,-0.0390625,-0.0078125,-0.078125,0,-0.03125,-0.0078125,-0.015625,-0.015625,-0.015625,-0.046875,-0.0078125,0.0078125,0.0625,0.0234375,0.015625,-0.03125,-0.015625,-0.046875,-0.0546875,0.03125,0.046875,-0.03125,0.015625,0.078125,0.046875,-0.03125,-0.0078125,0.0703125,0.0078125,0.015625,0.03125,0.0234375,-0.0078125,0.03125,-0.015625,0.0390625,-0.0234375,-0.0078125,0.015625,0,-0.0078125,0.0078125,0.0078125,0.0078125,0.015625,0,-0.015625,0.03125,0,-0.03125,0,-0.015625,0,-0.015625,0.046875,0.015625,0.046875,0,0.0234375,0.046875,-0.0546875,-0.046875,0.03125,-0.03125,-0.0390625,0.0078125,-0.0703125,0.03125,-0.046875,-0.0625,-0.0234375,0.0078125,0.0078125,0,0.0078125,0.0078125,0.0078125,0.0078125,-0.015625,0,0.03125,0.1015625,0.0390625,-0.03125,-0.0234375,0.0234375,-0.0078125,0,0,0,-0.0078125,0.0546875,-0.015625,0.0390625,0.015625,-0.0234375,-0.0078125,-0.0234375,-0.03125,0,0.0390625,-0.0078125,-0.0625,0.1015625,0,-0.0234375,-0.03125,0,0.046875,0,-0.0625,-0.03125,0.03125,-0.0078125,-0.0546875,-0.0234375,0.046875,-0.0703125,-0.015625,0.03125,0.0234375,0.0703125,-0.015625,-0.03125,0.03125,-0.03125,0.015625,0.046875,0.0078125,-0.0546875,-0.0078125,0.0078125,-0.0625,0,0.109375,-0.0390625,0,-0.0703125,-0.0078125,0.0078125,0.03125,-0.015625,-0.0078125,0.0390625,0,0.0390625,0.0703125,-0.046875,0.0078125,0,-0.0234375,-0.015625,0,0.0078125,0.03125,-0.015625,-0.0078125,-0.0390625,-0.0078125,-0.0390625,0.046875,0,-0.0703125,-0.03125,-0.0234375,-0.015625,-0.0234375,-0.046875,0,-0.03125,0.046875,0.015625,-0.09375,0.03125,-0.015625,-0.046875,0.0078125,0.046875,-0.03125,-0.078125,-0.0234375,0.0390625,0.0234375,-0.0234375,-0.03125,0.0390625,0,-0.015625,0.0234375,-0.0546875,0,0.0078125,-0.078125,-0.0234375,0.0859375,0.015625,0.0625,0,0,0.078125,-0.015625,-0.0546875,0,-0.015625,-0.0390625,-0.0234375,0.046875,0.0078125,-0.015625,-0.078125,-0.0390625,0.078125,-0.0234375,-0.046875,-0.015625,-0.0234375,0.0390625,0.0078125,0.0703125,0.0859375,0.0390625,-0.015625,-0.0546875,-0.0234375,0,-0.0078125,-0.0078125,0.0234375,-0.0078125,0,-0.015625,-0.0078125,0.0078125,-0.0078125,0.078125,-0.015625,0.078125,0.015625,0.046875,0.03125,-0.03125,-0.0625,-0.015625,-0.015625,-0.0234375,-0.0078125,-0.0078125,-0.078125,0.0078125,0.0390625,0.1953125,-0.0078125,-0.0703125,-0.046875,-0.015625,-0.046875,-0.046875,-0.0234375,0.078125,0.140625,-0.0078125,0.0078125,-0.0078125,0.0078125,0,0,0,0,0,-0.03125,-0.0859375,-0.1015625,-0.046875,-0.0625,0.0234375,0.03125,0.09375,0.0625,-0.0390625,-0.0625,0.046875,0,0.0546875,0.0234375,-0.015625,-0.0859375,-0.0078125,-0.03125,-0.0234375,-0.0234375,-0.1015625,0.0078125,-0.1484375,-0.0390625,-0.0078125,0.0234375,-0.0390625,-0.046875,-0.046875,-0.0078125,-0.0625,-0.0390625,0.0703125,-0.015625,0.0234375,-0.015625,-0.0625,-0.0234375,0.015625,0.0546875,-0.0078125,-0.0703125,0.0546875,0.03125,-0.015625,-0.0078125,0.0234375,0.0078125,-0.0234375,0.0625,0.0625,0.0703125,0.0390625,0.015625,0.015625,-0.015625,0.015625,0.0546875,0.0390625,-0.0390625,0.0078125,-0.0625,-0.015625,-0.03125,-0.0234375,-0.0390625,0,-0.0390625,0.0390625,0,-0.0078125,-0.03125,-0.015625,-0.0546875,0.0390625,-0.1171875,-0.078125,-0.0078125,0.15625,-0.046875,-0.0390625,-0.0234375,-0.03125,0.0625,-0.0859375,0.0703125,0.0234375,-0.0703125,-0.015625,-0.0078125,-0.0078125,0.0078125,0,-0.0078125,-0.015625,0.0078125,0,0,-0.0390625,-0.046875,-0.0078125,0.0234375,0.046875,-0.03125,0,-0.0390625,-0.0703125,0.046875,0.015625,0.015625,0,-0.046875,0.0234375,-0.0078125,-0.078125,0.09375,-0.0390625,-0.046875,-0.0234375,0.0546875,0,-0.0234375,0.03125,0.0234375,-0.015625,-0.03125,0,-0.0234375,0.0390625,-0.046875,0.109375,0.0234375,-0.0390625,0.0078125,0.0234375,-0.0390625,-0.0234375,-0.0625,-0.015625,0,0.03125,-0.03125,0.0390625,0.03125,0.0390625,0.0234375,0.078125,-0.09375,0.03125,0.0234375,-0.046875,0.0234375,-0.0078125,-0.0859375,-0.0234375,-0.1015625,0.0390625,-0.109375,0.0390625,0.0234375,0.0625,-0.046875,-0.03125,-0.015625,0.0703125,0.0859375,-0.0625,0.03125,0.0859375,0.0625,0,0.0625,0.0390625,-0.0390625,-0.015625,0.0078125,-0.09375,0.0078125,-0.140625,0.046875,-0.0078125,0,-0.0390625,0.03125,-0.03125,-0.03125,0.0078125,-0.0078125,-0.015625,-0.03125,-0.015625,-0.1484375,-0.0546875,-0.015625,-0.0234375,0.1015625,-0.1171875,0.0078125,-0.0078125,-0.03125,-0.046875,-0.1875,-0.015625,-0.0625,0.109375,-0.0546875,0.03125,-0.0390625,0.046875,-0.0234375,0.0078125,0.0078125,-0.078125,0.015625,-0.109375,-0.03125,0.0390625,-0.03125,0.0546875,-0.1015625,0.015625,0.0703125,0,-0.03125,0.015625,-0.0390625,0.046875,-0.0390625,0.0546875,-0.0625,0.0546875,0,-0.0390625,0.0390625,0.0703125,-0.015625,-0.0390625,-0.0703125,0,-0.015625,-0.015625,0,-0.0078125,0,-0.015625,-0.0078125,0.015625,-0.0078125,0,0.015625,0.0078125,-0.0234375,-0.109375,-0.1015625,-0.0078125,0.0234375,-0.0078125,0.0234375,-0.015625,0.0234375,0.046875,0.015625,0.0390625,-0.0390625,0.1015625,0.0078125,0.0234375,-0.046875,0.0625,-0.0078125,0.0390625,0.125,0,-0.109375,0.0078125,0.0390625,-0.03125,-0.0078125,-0.0078125,0.0078125,0,-0.0078125,0.0078125,0,0.0078125,0.0078125,-0.015625,-0.0703125,-0.015625,0.078125,-0.0546875,-0.0078125,0.0390625,0,-0.0625,-0.015625,-0.0078125,-0.0859375,-0.0234375,0.15625,0.0078125,0.078125,0.0390625,0.03125,0.03125,0.0234375,-0.1171875,0.0078125,-0.0078125,0.0078125,0.0390625,-0.0078125,-0.0078125,0.0078125,-0.0703125,-0.0703125,-0.0234375,0.03125,0.0234375,0,-0.0078125,0.03125,0.015625,-0.0625,0.0546875,0,0,-0.0390625,0.0234375,-0.0390625,0.015625,-0.0078125,-0.0078125,0.0078125,-0.0078125,-0.0390625,-0.015625,-0.0234375,0.015625,0.0078125,0.0234375,-0.015625,-0.015625,-0.0078125,0.0078125,0.03125,-0.015625,0.0078125,0.0078125,0.0234375,0.0234375,-0.0546875,0.046875,0.03125,0.03125,-0.09375,0.0078125,0.0078125,0.015625,0.0859375,-0.0078125,0.015625,-0.015625,0,0.03125,-0.09375,0.0078125,0.015625,-0.0234375,0.015625,-0.046875,0.0234375,0.078125,-0.0234375,0,-0.0078125,-0.015625,0,-0.0234375,0.0234375,0,0.0234375,0,0.0078125,0,-0.0078125,-0.0078125,0.015625,-0.046875,-0.0078125,0.0078125,-0.0234375,-0.015625,-0.0234375,-0.015625,0.0234375,0,0.0546875,0.0078125,-0.0390625,-0.0546875,0.0234375,0.0078125,0.015625,-0.0078125,-0.0625,-0.03125,0.015625,0.046875,0.046875,-0.0078125,-0.0390625,0.015625,-0.046875,-0.0234375,0.0234375,0.0078125,-0.015625,-0.0625,0.03125,-0.0390625,-0.015625,0.0234375,0.0234375,0.015625,0.015625,0.046875,-0.0390625,-0.0625,-0.0703125,-0.0078125,0.0078125,-0.0703125,0,0.0078125,-0.0546875,0.0234375,0.015625,-0.03125,-0.046875,0.0703125,-0.0078125,0.0703125,-0.0546875,-0.046875,-0.0546875,-0.03125,-0.0390625,0.0078125,-0.0390625,0.015625,0,-0.0234375,-0.015625,-0.015625,-0.0078125,-0.046875,-0.0390625,0.0390625,0.0390625,0.046875,-0.046875,-0.0234375,0.0546875,0.0078125,0.0234375,0,0.0078125,-0.03125,-0.015625,-0.0078125,0.078125,0.046875,0.0234375,-0.046875,0.0703125,0,-0.0234375,0.015625,-0.1171875,0.03125,-0.0625,-0.0234375,-0.0390625,-0.0546875,0,0.125,0.03125,0.078125,-0.0859375,0.0078125,0,0,0.0078125,0.046875,-0.1171875,0.03125,0.0390625,-0.015625,0.109375,-0.0234375,-0.0234375,-0.0078125,-0.078125,0.0234375,0.03125,0,-0.0234375,-0.015625,0.0390625,0.03125,-0.0078125,0.1171875,-0.078125,-0.015625,0.0703125,-0.0546875,-0.0703125,-0.015625,-0.015625,0.0234375,-0.0234375,0.0078125,-0.0390625,0.0625,-0.0546875,0.0625,-0.0703125,0.0078125,-0.03125,0,0,0,0.0078125,-0.015625,-0.015625,-0.0078125,-0.015625,-0.0234375,0.0078125,0.0625,0.0625,-0.0234375,0,-0.0546875,-0.0234375,0,-0.0078125,-0.0078125,-0.0078125,-0.0078125,-0.0078125,-0.046875,-0.0859375,0.046875,0.0078125,0.09375,0.0078125,-0.0625,0.109375,0.046875,0,-0.0546875,0,-0.0546875,0.078125,0.0078125,0.0234375,0.0078125,-0.0078125,0,0.0078125,0,-0.0078125,-0.015625,0.0703125,0.0703125,0.0390625,0.046875,-0.0859375,-0.0234375,0.09375,-0.0234375,0.03125,-0.0078125,0,-0.03125,-0.125,-0.078125,-0.078125,0.0234375,0,-0.0234375,0.0546875,-0.078125,0.015625,0.015625,-0.0703125,0.0078125,0.078125,-0.046875,0.0234375,-0.015625,0.0546875,-0.03125,0,-0.03125,0.03125,0.0078125,0.0625,0.015625,-0.0390625,0.0234375,-0.015625,0.0546875,-0.0234375,-0.0390625,0.0625,0,0.125,-0.0078125,-0.0078125,-0.0390625,0.046875,-0.0078125,-0.0078125,0.015625,-0.0390625,-0.046875,-0.0078125,-0.078125,-0.015625,0.0078125,0.046875,0.015625,0.0078125,0.015625,-0.0078125,0,0.0390625,-0.0234375,0.03125,-0.015625,-0.0078125,0.015625,0.0546875,-0.03125,0.0078125,-0.015625,0.0390625,0.046875,0.0390625,0.046875,-0.0078125,-0.0546875,-0.0078125,0,-0.03125,-0.0234375,-0.046875,0.1015625,-0.0234375,0.015625,0.0546875,-0.015625,-0.015625,-0.015625,-0.0078125,-0.03125,-0.0078125,-0.015625,0,0.0234375,-0.0078125,-0.015625,0.03125,0.015625,-0.0390625,0.0078125,-0.0078125,0,0,-0.0078125,-0.078125,0,0.0078125,-0.078125,0,0.046875,0.0234375,-0.0703125,-0.0078125,0.0234375,-0.0390625,-0.0078125,0.015625,0.0546875,0.046875,0.0234375,-0.09375,-0.046875,-0.0625,0.0234375,-0.03125,-0.046875,-0.03125,-0.0859375,-0.0078125,0,0,0.015625,-0.078125,-0.0078125,-0.0078125,-0.015625,0.0234375,0.0234375,0.046875,0.0859375,-0.0078125,0.0078125,-0.015625,0.0078125,-0.09375,0.03125,0.1015625,-0.046875,0.0234375,-0.078125,-0.09375,-0.046875,-0.0859375,0.0390625,-0.09375,0.15625,-0.0390625,0.0703125,-0.078125,0.0078125,-0.015625,0.046875,-0.0546875,-0.03125,0.0390625,-0.046875,0.0390625,-0.078125,-0.03125,-0.0234375,-0.03125,-0.0859375,-0.015625,0.0546875,0.0546875,0.0390625,0,0.03125,0.0390625,0,-0.0234375,-0.0390625,0.0078125,-0.015625,0,0.0859375,-0.0078125,-0.078125,-0.0703125,0.015625,-0.0703125,-0.015625,0.1484375,-0.0078125,-0.0390625,-0.03125,0,0.0390625,0.0546875,0,0,0,0.0078125,0.0234375,-0.0390625,-0.0078125,0,-0.1015625,-0.0625,0.234375,-0.046875,0.2109375,0.0078125,0.1171875,-0.0390625,-0.046875,-0.0234375,-0.015625,0.0078125,-0.1171875,0.0234375,-0.0546875,-0.046875,-0.109375,0.0703125,-0.0546875,0.03125,0.03125,0.0078125,-0.0546875,-0.0234375,-0.0390625,-0.046875,-0.015625,0.03125,0.03125,-0.015625,-0.0546875,-0.0390625,-0.0234375,-0.0078125,-0.0078125,0,0.0078125,-0.015625,0.0078125,0.015625,0.0078125,0.0234375,-0.046875,-0.0234375,0,0,0.015625,-0.015625,-0.0234375,-0.046875,0.0703125,0.03125,0.0234375,-0.015625,-0.0234375,-0.015625,-0.0078125,-0.03125,-0.0078125,-0.078125,0.109375,-0.0234375,-0.0234375,-0.0078125,-0.0234375,0.015625,0.0234375,-0.0078125,0.0078125,-0.0078125,0.015625,-0.0078125,-0.0078125,-0.0078125,0.0078125,-0.0078125,0,0.0703125,-0.046875,0,0.015625,-0.046875,-0.015625,0.015625,0,-0.046875,0.0390625,0.0078125,-0.015625,0.046875,-0.0234375,0.046875,-0.0078125,0.015625,0.0234375,0.09375,-0.0859375,-0.0390625,0.015625,-0.0234375,0.0078125,0.015625,-0.0390625,-0.0078125,0.046875,-0.0078125,-0.0078125,-0.0234375,-0.0546875,0,0,-0.03125,0,-0.015625,-0.015625,0.015625,-0.0078125,-0.0390625,-0.0625,0.046875,0.015625,0.03125,-0.0546875,0.0234375,0.015625,0.0078125,0.0078125,0.015625,0.015625,0.0078125,0,0.0078125,-0.015625,-0.03125,-0.0078125,0.0234375,0,0.0078125,0.0078125,0.0078125,-0.0078125,0.03125,-0.0078125,0.046875,-0.0078125,-0.0234375,-0.015625,0,0.015625,-0.015625,-0.0859375,0.0078125,-0.0390625,-0.0234375,0,-0.0234375,-0.0390625,-0.0234375,-0.0078125,-0.078125,-0.0625,0.0625,0.0078125,-0.015625,-0.0078125,-0.0078125,0,-0.0078125,-0.0078125,0.0078125,-0.015625,-0.0078125,-0.0078125,-0.0078125,0,0,0,-0.015625,-0.0234375,-0.015625,-0.0078125,0,0.015625,-0.0234375,0.0078125,0.0234375,0.0625,0.046875,-0.0078125,0.0078125,-0.0234375,0.0078125,-0.0546875,0,-0.0859375,-0.015625,-0.015625,0,0.0234375,0,-0.0234375,0.0078125,-0.0234375,-0.03125,-0.0078125,0.078125,0.015625,0.046875,-0.03125,0.0078125,0.03125,0.0234375,-0.0390625,0.0625,-0.03125,-0.015625,-0.0234375,-0.046875,-0.0234375,-0.0390625,-0.0234375,-0.078125,-0.0078125,0.0078125,0.03125,0.0078125,-0.0859375,-0.015625,-0.0234375,-0.0234375,-0.0546875,0.0859375,0.109375,0.03125,-0.03125,-0.0234375,-0.0546875,-0.0078125,0.0078125,-0.046875,0,-0.015625,-0.03125,0.0234375,-0.078125,0.0078125,0.0234375,-0.0234375,0.0078125,-0.015625,0.0234375,0.0234375,-0.0234375,0.046875,0.0234375,-0.0234375,0.015625,0.0234375,0.0390625,0.0078125,-0.0625,-0.0078125,0,-0.015625,0.03125,0.0078125,0.0234375,-0.046875,0.0625,0.015625,-0.0390625,0.0078125,-0.0078125,-0.0390625,0.03125,-0.03125,0.0078125,0.078125,-0.0234375,0,-0.09375,0.0078125,0.015625,0.015625,0.0703125,0.0234375,0,-0.015625,-0.046875,0.0078125,-0.046875,-0.0390625,-0.015625,-0.0078125,-0.015625,-0.0078125,0.03125,0.0390625,-0.0390625,-0.03125,0,-0.0078125,0.0078125,0.0859375,-0.0234375,0.0625,-0.0234375,-0.0390625,0.015625,-0.03125,0,-0.0234375,0.0234375,-0.0390625,-0.0390625,-0.015625,-0.0546875,0.0625,0.015625,-0.03125,-0.015625,-0.015625,-0.015625,-0.0078125,0,-0.015625,0,0.0078125,0.0078125,0,-0.09375,-0.0078125,-0.0390625,-0.09375,-0.015625,-0.015625,0.0546875,0,0.0390625,-0.0390625,-0.0078125,0.078125,-0.015625,0.0234375,0.0546875,-0.0390625,-0.0078125,-0.078125,-0.046875,-0.0625,0.0078125,-0.078125,-0.0234375,0.015625,-0.0703125,0.015625,0,-0.015625,0,-0.015625,0.015625,0,0,0,-0.0078125,-0.0078125,-0.09375,-0.0234375,0.046875,0,0.109375,0.015625,0,0.015625,-0.0078125,0.046875,-0.03125,-0.1015625,0.0078125,-0.0390625,0.03125,0.0625,0,-0.03125,-0.0546875,-0.0234375,-0.0703125,0,-0.015625,0.1171875,0.0859375,-0.046875,-0.0078125,-0.0703125,0.0078125,-0.0390625,0.03125,0,-0.03125,0.0390625,-0.0390625,-0.0078125,0.046875,-0.03125,0.046875,0.0078125,0.03125,0.0703125,-0.0390625,0.0234375,-0.015625,0.015625,0,-0.0546875,-0.0546875,-0.0390625,-0.0390625,-0.0078125,0.0234375,0.0234375,-0.03125,0.0078125,-0.0390625,0.0234375,-0.0390625,-0.0234375,-0.0078125,0.0078125,-0.015625,-0.0078125,-0.0234375,0.0390625,-0.0078125,0,0.0078125,0.0390625,-0.03125,-0.0234375,0.0703125,0.0390625,-0.0625,0.0546875,-0.0625,0.1171875,0.0078125,-0.0234375,0.0078125,-0.078125,0.046875,0.046875,-0.03125,0.0234375,0.0234375,0.0390625,0.0859375,0.015625,-0.0078125,-0.0078125,0.015625,0.0234375,0,0.0078125,0,-0.0078125,0.0546875,-0.0234375,0.0234375,-0.078125,-0.03125,-0.0078125,-0.0078125,-0.0234375,0.0078125,0.03125,0.0625,0,0.0625,0.0078125,-0.0546875,-0.015625,-0.0078125,-0.0234375,-0.046875,0.015625,-0.015625,-0.0078125,0.03125,-0.0703125,-0.046875,0.046875,-0.0390625,0.0078125,0.0234375,-0.03125,-0.03125,0.1640625,-0.0234375,-0.015625,0.0078125,-0.0390625,0,-0.03125,0.0390625,-0.015625,0.03125,0.0078125,0.03125,-0.078125,0.03125,0.0703125,-0.0078125,0.109375,0.0234375,-0.03125,0,-0.015625,0,-0.0078125,0.0234375,-0.015625,-0.0234375,-0.0859375,-0.0859375,-0.0703125,-0.015625,0.0390625,-0.0078125,0.0078125,-0.0390625,0.0078125,-0.0390625,-0.046875,-0.0703125,0.0078125,-0.0859375,-0.0078125,0.0390625,0.0234375,0.0234375,-0.0703125,0.0390625,-0.1015625,-0.0546875,0,-0.1015625,0.0234375,-0.0546875,-0.0078125,-0.03125,0.0390625,-0.0390625,-0.0078125,0.0078125,0.0234375,0.1328125,-0.140625,0.015625,0.0546875,-0.03125,0.0234375,-0.0234375,-0.125,-0.0234375,-0.0390625,-0.109375,-0.0859375,0.078125,-0.015625,-0.046875,0.078125,0.203125,0.03125,0.0234375,-0.1015625,-0.0625,0,0.03125,-0.015625,-0.0546875,0.0546875,0.0078125,0.0078125,0.03125,0.015625,-0.0546875,0,-0.03125,-0.0625,0.0703125,-0.0078125,0.1015625,-0.015625,0,0.0390625,0,0.03125,0,-0.0546875,0,0.0390625,0.03125,-0.0078125,-0.0078125,0.015625,-0.0078125,0,0.0234375,0,-0.0078125,-0.0078125,0.015625,0.0078125,0.015625,-0.0078125,-0.0078125,0,-0.0078125,0.1640625,0,0.015625,0.078125,-0.0546875,0.0078125,-0.0078125,0.0078125,0.03125,0,0.015625,0.0390625,0.015625,-0.0234375,-0.015625,-0.0078125,-0.0390625,0,0.0078125,-0.03125,0.0234375,0.0625,-0.015625,-0.0234375,-0.0625,-0.0234375,0.0078125,-0.015625,-0.0078125,0.0078125,-0.0078125,0.0078125,-0.015625,-0.015625,0.015625,0,0.0390625,0.0546875,0.0078125,0.0390625,-0.0390625,-0.0703125,-0.015625,0,-0.0078125,-0.0078125,0.015625,-0.0234375,-0.03125,0.0234375,-0.0390625,-0.03125,-0.03125,0.03125,0.0078125,-0.09375,0.015625,0.0546875,-0.015625,0.0078125,0,-0.015625,-0.0078125,0.015625,-0.015625,0.0078125,-0.03125,0.0078125,0,0.0078125,-0.0078125,-0.0078125,0,0.0625,-0.046875,-0.015625,0.09375,-0.0234375,-0.0390625,-0.0234375,0,-0.0078125,0.03125,-0.0078125,-0.0078125,0.0078125,-0.015625,0.015625,0.0390625,0,-0.03125,0,-0.0078125,-0.0390625,-0.0078125,-0.015625,-0.0078125,0,0.0234375,-0.015625,0.0078125,0.0078125,-0.03125,-0.046875,0.046875,0.0234375,0,0,-0.015625,0,-0.0390625,-0.0703125,0.0078125,-0.0078125,0,-0.0234375,0.0078125,0.078125,0.0234375,-0.0078125,-0.046875,0.0234375,0.0078125,-0.0078125,-0.046875,0.015625,0.015625,0.0390625,0,0,-0.0234375,-0.0078125,-0.015625,0.0078125,-0.015625,0.03125,-0.03125,-0.0078125,0.015625,0.015625,-0.03125,-0.0078125,0.015625,-0.015625,-0.015625,-0.046875,0.0078125,-0.0234375,0.015625,0.0078125,0.0234375,-0.0234375,-0.0078125,0.0703125,0,0.03125,-0.0859375,0.015625,-0.0546875,0,0,0.015625,0.0390625,0.09375,0.03125,-0.015625,-0.0625,-0.0078125,-0.0703125,-0.0546875,0.0234375,0.0703125,0.0859375,-0.046875,-0.0625,-0.03125,-0.0234375,-0.0625,-0.0546875,-0.03125,0.0234375,0.015625,-0.03125,0.015625,-0.0390625,0.0078125,-0.015625,-0.0078125,0,0.015625,-0.0625,-0.0078125,0.09375,-0.0625,0.0390625,-0.03125,-0.0390625,0.0234375,-0.0078125,-0.046875,-0.015625,0,-0.0234375,0.0078125,0.015625,0.015625,-0.0234375,-0.0859375,-0.015625,0.046875,-0.0390625,0,0.015625,0,0.0234375,0.015625,0.0703125,0.078125,0.0390625,0.0078125,-0.046875,-0.0078125,-0.0234375,-0.0234375,0,-0.1015625,-0.0234375,-0.015625,-0.0625,-0.0234375,0.0390625,-0.0078125,0.046875,0.015625,0.03125,0.03125,0.0078125,0,-0.0546875,0.0078125,-0.0390625,-0.03125,0.015625,0.046875,0.0234375,0.015625,0.03125,-0.0078125,0.0078125,0.0390625,-0.0625,-0.0234375,0.0859375,0,0.015625,0.0078125,-0.03125,-0.015625,-0.015625,-0.015625,0,-0.0234375,0.03125,-0.0390625,-0.078125,0.0234375,0,-0.03125,-0.03125,0,0.046875,0.0546875,-0.03125,-0.078125,0.09375,-0.0859375,0.0078125,-0.0234375,0.046875,0.0078125,0,0.015625,0.0078125,0,-0.0234375,-0.015625,0.0078125,0,-0.0234375,0,0,-0.0078125,0.015625,0.0234375,0,-0.03125,0.015625,-0.03125,-0.0078125,0.0546875,0.03125,-0.015625,-0.03125,0.0234375,-0.0234375,-0.015625,-0.0625,-0.0078125,-0.046875,0.015625,0.0234375,-0.015625,-0.015625,-0.03125,-0.0078125,0,-0.015625,0,0.0078125,0.0078125,-0.0078125,0.0078125,-0.0078125,0,-0.0234375,-0.015625,-0.015625,0.0703125,-0.09375,-0.1015625,0.015625,-0.0234375,-0.0546875,0.0546875,0.0078125,0.0390625,-0.0546875,0.0078125,-0.015625,0.046875,-0.0078125,0.0234375,0.0234375,0.0234375,-0.03125,-0.0390625,-0.078125,-0.046875,-0.0859375,0,0.046875,0.015625,-0.125,-0.046875,-0.0546875,0.03125,0.1015625,-0.046875,-0.0234375,0.0546875,-0.0234375,-0.0078125,-0.0234375,0.0390625,0.0078125,0.0546875,0.0703125,0,0.0625,0.0390625,0.0234375,-0.015625,-0.03125,-0.0234375,-0.03125,-0.046875,-0.015625,-0.0078125,0.0234375,0.0390625,0.046875,-0.0078125,-0.0078125,0.015625,-0.015625,0,-0.015625,-0.015625,0.0390625,0.03125,-0.0234375,-0.015625,-0.0234375,0,0.09375,-0.0390625,0.078125,-0.03125,0.0390625,-0.0234375,-0.046875,-0.0234375,0.015625,0.0234375,0.1015625,0.0078125,-0.046875,-0.1015625,0.0625,-0.0390625,0.015625,-0.03125,-0.0234375,0.0390625,0,-0.015625,-0.0078125,0.0234375,0.0234375,0.0234375,0.0234375,0.0078125,0.0234375,0.015625,-0.0234375,-0.0078125,-0.0234375,-0.015625,-0.015625,0.0078125,-0.0078125,-0.0234375,0.0234375,0,0.1171875,0.0390625,-0.0546875,-0.046875,0.0390625,0.0390625,0.03125,0,0.0078125,0.0234375,-0.078125,0,0.015625,-0.0703125,-0.0625,-0.046875,0.046875,-0.09375,0.046875,-0.0078125,0.0234375,0.0390625,-0.0546875,0.0234375,0.015625,0.0390625,0.03125,0.0078125,-0.0234375,-0.0390625,-0.015625,0.0546875,-0.125,0,0.0390625,0.0234375,0.0703125,-0.0234375,-0.0078125,-0.046875,-0.0078125,0.0234375,0.0234375,0.0625,0.0546875,0.046875,-0.03125,-0.0703125,-0.0078125,-0.0390625,0.015625,-0.0234375,-0.0078125,0.0234375,0.015625,-0.0625,0.03125,-0.0078125,0.0078125,-0.0625,0.046875,0.0390625,0.0234375,0.0703125,-0.0078125,0.046875,-0.0703125,0.0234375,-0.015625,0.09375,0.046875,0.046875,0.0859375,-0.0078125,-0.0234375,-0.015625,0.0234375,0.0625,-0.078125,-0.03125,-0.0703125,0.015625,0.0546875,-0.078125,0.0625,0.0078125,0.03125,0.03125,-0.0078125,-0.0546875,-0.046875,-0.0078125,-0.0546875,0.03125,0.0234375,0.1015625,0.0703125,0.03125,0,0.03125,-0.0234375,0.03125,0.0703125,-0.0078125,0.03125,0.015625,-0.03125,-0.0078125,0.046875,-0.0625,0.0390625,-0.0078125,0,0.0234375,-0.0234375,0.0625,0.0546875,0.0703125,0.0078125,-0.0546875,-0.0546875,-0.09375,-0.1171875,-0.046875,0,0.015625,0.0078125,0.0078125,-0.03125,0.015625,-0.015625,0.046875,0.0859375,0.015625,-0.0078125,0.0078125,-0.0078125,-0.0078125,0.0234375,0,0.0078125,-0.0078125,0,-0.0078125,0.015625,0.0078125,0.015625,-0.03125,-0.0859375,0,-0.0234375,0.0078125,-0.0078125,0.015625,0.09375,-0.046875,0.0546875,0,-0.015625,0.0234375,-0.0078125,0.0234375,0,-0.0078125,0.0390625,-0.015625,-0.015625,-0.0625,-0.03125,-0.0078125,-0.0078125,0.0078125,-0.015625,-0.015625,-0.015625,0,0,0.0078125,-0.0234375,-0.0234375,-0.0234375,0.0078125,-0.09375,-0.046875,0.1015625,-0.0703125,0.0078125,-0.0078125,-0.0390625,-0.0078125,-0.1015625,0,0,0.1171875,0.0703125,0.0703125,-0.015625,-0.0234375,0,0.0078125,-0.0234375,0.0078125,-0.015625,-0.0546875,-0.03125,0.0078125,-0.0078125,-0.03125,-0.0234375,0.0625,0.015625,0.0078125,0.0390625,0.03125,0.0078125,-0.046875,0.0078125,0.0234375,-0.015625,-0.0234375,-0.0390625,-0.015625,0.03125,-0.015625,-0.0234375,-0.0078125,0.015625,0.0078125,0,-0.015625,-0.0234375,-0.0078125,-0.0078125,-0.0234375,-0.0078125,0.0078125,-0.0390625,0.015625,0.0234375,-0.015625,0.0078125,0.0390625,0.015625,-0.0078125,-0.0078125,0.046875,0,-0.0234375,0.0234375,-0.0234375,0.03125,0.015625,0.0078125,-0.0703125,-0.0390625,-0.09375,0.171875,-0.1171875,0.0234375,-0.03125,-0.0078125,-0.015625,-0.0546875,-0.0546875,0,0.0546875,-0.109375,0.0625,0.015625,0.0234375,-0.0078125,-0.0078125,0.0078125,0,0,0.0078125,0,0,-0.0078125,-0.0078125,0.015625,0.015625,-0.0078125,0.015625,0.0234375,-0.0234375,0.0234375,-0.0234375,-0.0234375,-0.03125,-0.0859375,0.015625,0.0390625,0.0390625,0.046875,-0.0234375,-0.0234375,-0.03125,-0.0703125,0.0078125,0.0078125,-0.03125,0,0.0078125,0.03125,0,-0.0546875,-0.140625,0.03125,-0.03125,-0.015625,0.0546875,0.0234375,-0.015625,-0.046875,-0.0390625,-0.0078125,-0.09375,-0.0078125,0.078125,-0.0234375,0.09375,-0.03125,-0.0234375,0.0078125,-0.015625,-0.0546875,0.078125,0,-0.0390625,-0.0390625,-0.03125,-0.0078125,-0.015625,0.0546875,0.0078125,0.0390625,-0.0390625,-0.0625,-0.0234375,-0.0234375,0,-0.015625,-0.0078125,0,-0.015625,-0.0546875,-0.046875,-0.0546875,0.0390625,0.0546875,0.015625,-0.015625,0.015625,-0.03125,0.03125,-0.0078125,0.0390625,-0.0078125,0.015625,0,0.0390625,0.0234375,0.09375,-0.0390625,0.0234375,0.0234375,0,-0.03125,-0.0234375,0.0546875,-0.1015625,0.09375,0.046875,-0.046875,0,0.0234375,0,-0.046875,-0.0703125,0.046875,-0.0078125,0.09375,0.03125,0.03125,0.0078125,-0.0234375,0,0.078125,0.015625,0.0234375,-0.0625,-0.0390625,-0.015625,-0.0234375,-0.03125,-0.0078125,-0.0390625,0.1640625,-0.03125,0.03125,0.0078125,-0.03125,-0.0703125,-0.0234375,-0.0234375,0.1171875,-0.0625,0.046875,-0.0625,-0.0703125,-0.0078125,-0.046875,0,0,-0.0390625,-0.015625,-0.0078125,-0.0234375,-0.0078125,0.0078125,0.015625,-0.0078125,-0.0078125,0.0234375,0.015625,-0.015625,-0.0078125,-0.0078125,0,-0.0078125,0.015625,0.0078125,0.0234375,-0.0234375,-0.0234375,0.03125,-0.015625,-0.0078125,-0.0234375,0.0546875,-0.0078125,-0.0078125,0.015625,0,-0.015625,0.015625,0,-0.0546875,0.0390625,-0.0078125,0,0.0078125,-0.015625,0.03125,0.0390625,-0.0234375,-0.0078125,0,0.0078125,0.015625,-0.0078125,0.0078125,-0.0078125,-0.0078125,0,-0.0390625,0.0546875,-0.015625,-0.03125,0.0390625,-0.015625,0.078125,0.03125,0,0.0390625,-0.046875,-0.0078125,0.03125,-0.0546875,-0.0234375,-0.046875,-0.0234375,-0.0078125,0.03125,0,-0.0078125,-0.09375,0,0,0.015625,-0.015625,-0.0078125,0.046875,-0.0234375,-0.0078125,0.0390625,0,-0.0234375,0.046875,0.015625,0,0.015625,-0.0390625,-0.015625,-0.0234375,-0.015625,0,0.0234375,-0.03125,0.015625,-0.0625,-0.046875,0.0078125,0,-0.0390625,0,0.0078125,-0.0078125,-0.015625,-0.015625,-0.0234375,0,-0.0078125,0,-0.0078125,0,0.0078125,-0.015625,-0.03125,-0.0078125,0,-0.03125,0.015625,-0.015625,0.03125,-0.03125,0,-0.0546875,-0.0546875,0,0.078125,0.0078125,0.015625,-0.0625,-0.015625,-0.015625,0.046875,0.09375,-0.015625,-0.1015625,0.0390625,-0.015625,0.0078125,0.0390625,-0.015625,0.015625,0.0078125,-0.015625,-0.0078125,0,0,0,-0.0078125,-0.0078125,-0.03125,-0.0546875,0.0078125,0.0078125,0.015625,-0.0078125,0.0078125,-0.0078125,0.0078125,0,-0.0234375,0,0.0390625,-0.0859375,0,0.0625,0.0234375,-0.0078125,0.0703125,-0.046875,0,0.1484375,-0.078125,-0.0078125,-0.0234375,0.0078125,0,-0.0546875,0.0078125,-0.015625,-0.015625,0.0078125,-0.03125,-0.046875,0.046875,0,-0.0234375,-0.0234375,-0.0078125,-0.0546875,0.0390625,-0.0234375,0.0390625,0.0625,-0.0234375,-0.0546875,-0.0234375,-0.0078125,-0.0625,-0.03125,-0.0078125,-0.0390625,0.0234375,-0.0078125,-0.078125,-0.0078125,0,0.078125,-0.0546875,-0.015625,-0.0234375,-0.0234375,0.0078125,0.03125,-0.0078125,0,-0.0234375,0.046875,-0.0234375,-0.0390625,-0.015625,0,-0.03125,-0.0078125,0.0078125,-0.015625,-0.0234375,0,-0.0234375,0.0078125,-0.015625,-0.015625,-0.0078125,-0.0078125,-0.03125,0.0078125,-0.015625,0.0390625,-0.0078125,-0.0078125,-0.015625,-0.0625,0.015625,-0.03125,0.015625,-0.0234375,0,-0.0546875,-0.0234375,0.015625,0.0859375,0,0.09375,-0.0234375,-0.03125,-0.0625,-0.0078125,-0.0234375,-0.046875,0.0625,-0.0078125,0.015625,-0.015625,-0.0234375,0.015625,-0.078125,0,0.015625,0,-0.0078125,0.046875,-0.0234375,-0.0078125,-0.015625,0.0234375,-0.0078125,-0.0625,-0.0546875,0.015625,0.0078125,-0.078125,-0.0234375,0,0.015625,-0.015625,-0.0234375,-0.015625,-0.0234375,0.03125,0.015625,0.046875,0.0078125,0.046875,-0.0390625,-0.0078125,-0.015625,0.0078125,-0.0078125,-0.0078125,-0.0078125,0,0.0078125,0,-0.015625,-0.046875,0.078125,0.0625,-0.0390625,-0.015625,-0.0390625,0.0078125,-0.0546875,-0.0078125,-0.015625,-0.015625,0,0.015625,-0.015625,-0.0546875,-0.0390625,-0.015625,-0.0078125,0.0078125,0.015625,0.0859375,-0.0078125,-0.03125,-0.0234375,0,-0.0234375,-0.0078125,0.0078125,0.0078125,-0.0078125,-0.015625,0.015625,0.0078125,-0.0078125,0.0078125,-0.0390625,0.0078125,-0.0234375,-0.015625,-0.0234375,-0.078125,-0.015625,-0.0546875,0,0.0625,0.109375,-0.0078125,0,0.0390625,-0.0546875,-0.0234375,0.0078125,0.0078125,-0.0234375,0.0234375,-0.0078125,0,-0.046875,-0.015625,-0.0546875,-0.046875,-0.0078125,0.0078125,0.015625,0.0078125,0,0.0234375,-0.0390625,-0.0078125,0.0390625,-0.0234375,0.0234375,0.0703125,0.0390625,-0.0546875,-0.03125,-0.0390625,0.03125,0.046875,-0.0234375,0,0.03125,-0.0234375,0.015625,0.015625,-0.0234375,-0.015625,0.0078125,-0.0234375,-0.046875,0.0390625,0.0078125,-0.015625,0.015625,0.015625,0.0078125,0.015625,0.0078125,-0.0078125,0,0,-0.0078125,-0.0390625,0.0078125,0.0234375,-0.0390625,0.0078125,-0.0390625,-0.0234375,0.0078125,-0.015625,-0.0234375,0.0234375,-0.015625,0.03125,-0.046875,-0.0546875,-0.0390625,0.0078125,-0.0234375,-0.0546875,0.0546875,0.015625,0.015625,-0.03125,0.0078125,0.0078125,0.0078125,0.0234375,0.015625,0.0078125,0,0,0,0.0078125,-0.015625,-0.0078125,-0.015625,0,-0.0390625,-0.0078125,0,0,-0.0078125,-0.015625,-0.0234375,-0.015625,-0.0234375,0.0078125,0.0703125,-0.0234375,0.0234375,0.015625,0.0078125,0,-0.015625,-0.0703125,0.0234375,-0.0390625,-0.0234375,-0.015625,0,0.015625,-0.0234375,-0.0625,-0.109375,0.015625,0.109375,0.03125,-0.0078125,-0.015625,0.0234375,-0.0390625,-0.0234375,-0.0078125,0,-0.0234375,0.0625,0.0078125,-0.046875,-0.0234375,0.0234375,0.0625,0.0859375,0.0234375,-0.0078125,-0.03125,0,-0.015625,0.0078125,-0.03125,-0.015625,-0.03125,0.015625,0.046875,-0.109375,0.078125,-0.0546875,-0.015625,0,-0.0234375,-0.0625,-0.0078125,0.0078125,0.03125,0.0078125,0.0234375,-0.03125,0.03125,0.0546875,-0.0390625,-0.015625,-0.0390625,-0.0078125,0.03125,0.03125,0.0703125,-0.0390625,0.0234375,-0.03125,0.015625,0,-0.0390625,0.0234375,-0.0234375,-0.0703125,0.015625,-0.046875,-0.0390625,-0.046875,0.0703125,0.0390625,-0.0546875,0.03125,0.03125,0.046875,0.046875,0.0078125,-0.03125,0.046875,0.0234375,-0.0703125,0.0078125,0.03125,0.0625,-0.015625,0.015625,-0.0234375,-0.03125,-0.03125,0.0234375,0.0078125,-0.015625,0.0078125,0.0390625,-0.0390625,-0.0078125,-0.0390625,-0.0390625,0,0.0078125,0.015625,-0.0390625,-0.03125,0.015625,-0.046875,-0.015625,-0.0078125,0.015625,-0.0546875,-0.0078125,-0.015625,-0.0078125,0,0.015625,0.0078125,0.0625,-0.0078125,-0.0078125,0.0078125,-0.0078125,0,0.0078125,0,0,-0.015625,0.0078125,-0.015625,-0.0703125,0.0234375,-0.03125,0.0078125,-0.0234375,0,0.0234375,0.0390625,0.0234375,-0.03125,0.03125,-0.0390625,-0.078125,-0.0078125,0.046875,0.015625,0,0.0078125,0.03125,0.0234375,-0.0703125,0.015625,-0.0546875,0.0390625,-0.0078125,0.0234375,-0.0078125,-0.0078125,-0.015625,-0.0078125,0,0.0078125,0.0078125,-0.015625,0.0078125,0,-0.0234375,0.03125,-0.015625,0,0.0078125,0.0546875,0.015625,0.0234375,-0.078125,-0.0078125,-0.046875,0.0546875,-0.078125,-0.0078125,-0.0078125,-0.03125,0.0703125,-0.0625,0.046875,-0.0234375,-0.0234375,0.015625,-0.0546875,-0.046875,0.09375,-0.0078125,-0.03125,-0.015625,-0.046875,-0.03125,0.0546875,0.015625,-0.0703125,-0.0390625,-0.0390625,0.0390625,0.03125,0.0390625,0.015625,-0.0234375,-0.0390625,-0.046875,0.03125,0.0390625,-0.015625,-0.015625,-0.03125,0.03125,-0.0078125,-0.0390625,0.0546875,0.0078125,0.03125,-0.046875,-0.046875,-0.0078125,0.0390625,0.0078125,-0.015625,0.046875,-0.0078125,0,-0.0078125,-0.0078125,0.03125,-0.0234375,-0.0078125,0.03125,0,0.078125,-0.0078125,-0.0078125,0.0390625,0.0078125,-0.03125,-0.1015625,0.03125,0.0546875,-0.03125,0.0703125,0.0390625,-0.0390625,0.0078125,-0.015625,-0.0703125,0.03125,-0.109375,-0.03125,-0.0546875,0.0078125,0.0234375,0.0078125,0.0078125,0.0234375,0.03125,0,0,0.0078125,0.015625,0.0078125,-0.0078125,0.015625,0.078125,-0.0078125,0.0078125,0.0546875,0.0078125,0.046875,0.03125,0.0859375,0.0234375,-0.0546875,-0.0234375,0.0625,-0.046875,-0.0078125,0.015625,-0.015625,0.0078125,-0.046875,-0.1015625,0,0.0625,0.09375,0.0390625,-0.0234375,0.015625,0.0390625,0.0234375,-0.0625,-0.046875,0.1015625,0.015625,0.0859375,-0.03125,-0.03125,0.0078125,-0.0234375,-0.0078125,0.0234375,-0.0625,0,-0.0390625,0.015625,-0.03125,0.0390625,-0.015625,0.0625,-0.0703125,0.0546875,0.0078125,-0.0546875,0.03125,-0.0703125,0.0625,0.0625,-0.109375,-0.0078125,0.015625,-0.0546875,0.0234375,-0.0078125,0.09375,0.03125,-0.0546875,0.09375,0,-0.015625,0.0390625,-0.0078125,-0.046875,0.015625,0.0546875,0.0390625,-0.0078125,-0.046875,0.0546875,0.015625,0.046875,-0.03125,-0.0703125,0.03125,0.0234375,-0.0546875,-0.0390625,-0.0703125,-0.03125,0,0,0,0.09375,-0.046875,-0.015625,-0.0703125,-0.015625,0.0234375,-0.0234375,0.0390625,0.015625,0.0234375,0.0390625,-0.078125,-0.0390625,0.109375,-0.0703125,0.09375,0.0078125,-0.0625,0.046875,0.03125,-0.0859375,-0.0546875,-0.03125,-0.015625,-0.0390625,-0.015625,-0.0859375,-0.0234375,0.1171875,-0.0625,-0.046875,0.015625,-0.046875,0,0.0234375,-0.0234375,0.0234375,0.0234375,-0.0625,-0.03125,-0.0703125,-0.0078125,0,-0.0234375,-0.015625,0,0.0546875,0.046875,0.0234375,-0.09375,-0.0703125,0.015625,0.0078125,0,0.0078125,-0.0078125,0,-0.0078125,-0.0078125,-0.015625,0,-0.015625,-0.015625,-0.0390625,0.046875,-0.0234375,-0.0234375,0.0625,0,-0.0078125,-0.0390625,0.015625,0.0078125,0.046875,-0.0234375,0.046875,0.046875,-0.015625,0.0078125,0.0234375,0.0546875,0.03125,0.0078125,-0.0703125,0.015625,-0.015625,-0.0078125,-0.03125,-0.0078125,-0.0078125,-0.0078125,-0.0078125,0,0.0078125,-0.015625,-0.0078125,0.0078125,-0.0234375,-0.0078125,-0.015625,0.0390625,0.0234375,0.0546875,0.046875,-0.015625,-0.0078125,-0.0078125,0.078125,0.0546875,-0.0390625,0,0.0390625,-0.015625,0.0078125,-0.0078125,-0.0078125,0.046875,0.015625,-0.046875,-0.015625,-0.0390625,0.0390625,-0.015625,-0.0234375,0.015625,-0.0390625,-0.0625,0.0078125,0.015625,-0.0234375,-0.046875,-0.0546875,-0.03125,-0.0078125,0.0078125,0.015625,0.078125,-0.03125,0.046875,-0.078125,-0.0078125,0.015625,0.015625,0,0.0234375,-0.046875,0.0703125,0.015625,-0.0078125,0.0078125,0.015625,0.0078125,0,0,-0.03125,0.03125,-0.03125,0.0078125,0,0.0078125,-0.0234375,0.0390625,-0.0234375,-0.078125,-0.03125,-0.0234375,0.0078125,0.03125,0.015625,-0.0546875,-0.0234375,-0.046875,0.0859375,0.0546875,0.0078125,-0.0390625,-0.0625,0.0078125,0.015625,-0.0234375,-0.015625,0.1328125,-0.015625,-0.09375,0.0625,-0.0078125,0.0078125,0,0,0.015625,0.03125,-0.015625,0.015625,0.0234375,-0.0078125,0,-0.0390625,-0.015625,-0.0234375,0.0078125,-0.015625,0.0234375,0.0234375,0.0078125,-0.015625,-0.03125,-0.0078125,-0.015625,0.0546875,0,-0.03125,0.0234375,-0.0078125,-0.046875,0.015625,-0.0234375,-0.03125,-0.0546875,0.03125,-0.03125,0.0234375,0.015625,-0.015625,-0.0390625,-0.046875,-0.015625,0.03125,-0.0234375,-0.0234375,0.0703125,0.078125,0.03125,0.046875,-0.046875,0,-0.0234375,0.03125,-0.0078125,0.015625,-0.046875,-0.046875,0.0078125,0,-0.0078125,0.1328125,-0.0234375,0.0546875,0.09375,0,0,-0.0234375,0,0.015625,-0.0390625,-0.0625,-0.0625,0.1328125,0.0859375,-0.046875,-0.0390625,-0.0625,0.03125,-0.0625,-0.0703125,-0.0234375,0.0078125,0.015625,0.0078125,0.078125,0.078125,0.015625,-0.0234375,0.0234375,0.015625,-0.0078125,-0.0390625,-0.0390625,0.046875,0,0.015625,-0.0078125,0.109375,-0.0546875,0,-0.0078125,-0.015625,-0.0234375,0.078125,0.0234375,-0.109375,-0.015625,-0.0390625,0.0546875,-0.015625,-0.0078125,-0.0078125,0.0546875,-0.0390625,-0.0078125,-0.0625,-0.046875,-0.0546875,-0.0390625,-0.03125,0.078125,-0.0234375,0,0.0078125,-0.0703125,0.015625,0.015625,0.0078125,-0.046875,0.046875,-0.0625,-0.0546875,0,-0.0234375,-0.03125,0.0078125,0.015625,0.0078125,-0.0625,-0.0234375,0.015625,-0.0625,-0.0625,-0.015625,0.0078125,0,-0.0390625,0,0.0390625,0.0703125,-0.015625,0.0703125,-0.03125,-0.015625,-0.0078125,-0.0703125,0.0078125,0,-0.0078125,0.0078125,0.015625,0.0078125,0.015625,0,0.015625,0,0,-0.0234375,-0.03125,-0.109375,-0.09375,0.0234375,0.015625,0.109375,-0.03125,0.03125,0,-0.0546875,-0.0390625,0.0078125,-0.0546875,0.046875,0.0234375,0.015625,0,0.0078125,-0.015625,0.0234375,-0.0703125,-0.0390625,-0.0078125,0.0234375,-0.0078125,0,-0.0078125,0.0078125,-0.0078125,0.0234375,0,0.0078125,-0.0078125,0,-0.0546875,-0.0234375,-0.0703125,-0.0234375,-0.0546875,-0.015625,0.15625,-0.0390625,0,0.0234375,-0.0703125,-0.0078125,-0.1796875,0.15625,-0.0078125,-0.1015625,0.0546875,0.0078125,-0.0234375,0.0625,0.0078125,0.0234375,0.03125,-0.0625,0.0234375,-0.0859375,0.015625,0.015625,-0.0078125,-0.0078125,-0.0859375,0.0390625,0.0078125,-0.015625,-0.0234375,-0.015625,-0.0546875,0.0234375,-0.0234375,0.0859375,0.046875,0.03125,0.1171875,-0.078125,0.015625,0,-0.03125,-0.03125,0.0078125,0.0078125,0.015625,-0.03125,0,-0.0234375,0.0234375,0.046875,0.0078125,-0.03125,0,-0.0078125,-0.0234375,-0.0078125,0.015625,0.0078125,-0.046875,0.0078125,-0.0234375,0,0.0234375,0.046875,0.0859375,-0.0078125,-0.03125,0.0234375,-0.0546875,0.0078125,-0.09375,-0.015625,0.0234375,0.0859375,-0.0234375,0,0.1015625,-0.0234375,-0.03125,-0.0234375,-0.046875,-0.015625,-0.1015625,-0.0078125,0.0078125,0,-0.0078125,0,0,0,-0.0078125,-0.03125,-0.0078125,0.0234375,-0.0390625,0.0078125,-0.0078125,-0.0078125,0.0078125,0,0.03125,-0.0078125,0.0390625,-0.03125,-0.0234375,0.046875,0.03125,-0.0703125,0.0078125,-0.0078125,-0.0078125,-0.078125,-0.078125,-0.046875,0.0390625,0.0234375,-0.03125,-0.09375,0.2109375,0.0390625,0.0703125,0.0546875,0,-0.0078125,-0.0703125,-0.015625,-0.0078125,0.046875,-0.03125,0.015625,0.015625,-0.0390625,-0.046875,-0.0859375,0.015625,0.03125,-0.0390625,-0.0078125,0.03125,0.0703125,-0.0390625,0.0078125,-0.0546875,-0.03125,-0.03125,-0.015625,-0.0390625,0.0703125,-0.1015625,-0.046875,0.0390625,0.0234375,-0.0234375,-0.09375,0.109375,0.0078125,-0.03125,0.0078125,-0.0078125,0.0546875,0.0625,-0.03125,0.015625,-0.046875,-0.0234375,-0.0078125,0.0234375,0.015625,-0.03125,-0.0078125,-0.015625,-0.0234375,-0.015625,-0.0546875,-0.0625,-0.1171875,-0.0625,-0.03125,0.0625,-0.0234375,0.0078125,0.0625,0.0625,0.0546875,-0.015625,-0.0234375,-0.109375,-0.03125,-0.0234375,0.0546875,-0.0234375,0.0234375,0.078125,-0.0234375,-0.0390625,-0.03125,-0.0234375,-0.03125,0.015625,0.0703125,-0.0234375,-0.046875,-0.0078125,0.015625,-0.03125,-0.03125,0.0390625,-0.0625,0.03125,-0.0078125,0.03125,0.0546875,0,0,0,-0.03125,-0.0234375,0.046875,0,-0.015625,-0.078125,-0.015625,-0.046875,0.09375,-0.03125,-0.046875,0.0234375,-0.0390625,-0.015625,-0.0234375,0.015625,-0.015625,-0.03125,0.046875,-0.0234375,0.03125,-0.015625,-0.015625,-0.015625,-0.015625,-0.015625,-0.0078125,0.015625,0.0078125,0.0078125,-0.015625,0.0078125,-0.046875,-0.0234375,-0.0546875,0,0.078125,0.046875,-0.015625,0.015625,0.015625,-0.046875,0.0078125,-0.015625,0.015625,0.015625,0.0859375,-0.0078125,-0.0234375,-0.0078125,0,0,-0.0546875,0.0078125,0.078125,-0.0546875,0.09375,0,0.0078125,0.0078125,-0.0078125,0,0.0078125,0,0.0078125,0,-0.0078125,0.015625,0.03125,-0.0390625,-0.0546875,0.0234375,-0.0390625,0.1328125,-0.046875,-0.0546875,0.03125,-0.03125,-0.09375,0.0859375,0.0078125,-0.0546875,0.03125,0.09375,0.078125,-0.03125,0.0078125,0.0859375,-0.109375,-0.0078125,0.0234375,0,-0.0546875,0.0546875,-0.0234375,0.0234375,-0.0390625,0.015625,-0.0234375,0.0078125,0.0234375,-0.0234375,0.03125,-0.0234375,-0.015625,0.0234375,-0.0546875,0.015625,-0.0234375,-0.015625,0.0078125,-0.015625,-0.015625,0.03125,-0.015625,0.03125,-0.0390625,0,-0.0078125,0.03125,-0.03125,-0.046875,0.015625,0.0078125,0,0.0078125,0.015625,-0.0078125,-0.015625,0.0546875,0.046875,-0.0078125,0.0234375,0,-0.0234375,0.015625,-0.0078125,-0.015625,0.015625,0.0078125,0.015625,0.0390625,-0.0625,-0.0390625,-0.0078125,0.09375,0.0078125,-0.015625,-0.0078125,-0.0078125,0.0390625,-0.03125,-0.078125,0.0078125,0.015625,-0.046875,-0.0078125,0,-0.0078125,-0.0078125,-0.0078125,0.015625,-0.0078125,-0.0078125,-0.015625,0.015625,0.015625,0.015625,-0.0078125,0.015625,0.015625,-0.0234375,0.0625,0,0.0390625,0.0078125,0,-0.0234375,-0.0234375,0,-0.03125,-0.046875,0.03125,-0.03125,0,0.0078125,-0.015625,-0.0546875,-0.0078125,-0.0078125,-0.015625,-0.046875,0.0078125,-0.0546875,-0.046875,-0.03125,-0.0625,0.0078125,-0.046875,-0.0859375,0.046875,-0.015625,-0.0234375,0.0625,-0.0078125,0.03125,-0.03125,0.0703125,-0.078125,0.0234375,0.015625,0.046875,-0.03125,0.03125,-0.0390625,-0.0078125,-0.0078125,0.046875,-0.015625,0.1015625,0,-0.0078125,-0.046875,-0.03125,0.015625,0.0234375,-0.03125,0.0234375,0.015625,0.0390625,0.0546875,-0.0390625,-0.0078125,-0.0078125,0.015625,0.03125,0.0390625,0.0546875,0.0234375,-0.0078125,0.03125,-0.0390625,0.0234375,-0.0234375,-0.015625,0.0390625,0.0234375,-0.03125,-0.0390625,0.0390625,0.0234375,-0.0234375,0,-0.03125,-0.0234375,0.109375,0.0234375,0.0390625,-0.0234375,-0.0546875,-0.0390625,-0.0625,-0.015625,-0.015625,0.0234375,-0.0234375,-0.03125,-0.0703125,-0.015625,-0.046875,0.0390625,-0.0078125,0.0546875,-0.015625,0.015625,-0.0546875,0.046875,0.0078125,0,0.015625,0.0546875,0.0390625,-0.0546875,0.0078125,-0.078125,-0.03125,-0.0625,0,-0.0078125,0.046875,0.0078125,0.015625,0.046875,-0.015625,0.0078125,-0.046875,0,0,-0.0234375,0.0859375,0.0234375,0,0,-0.046875,-0.046875,-0.0234375,0,-0.0078125,-0.015625,0.0078125,-0.0078125,0.0078125,0.0078125,-0.015625,-0.015625,-0.015625,-0.0078125,0.015625,-0.046875,-0.0234375,-0.046875,0.0390625,0.0390625,-0.0234375,-0.0625,-0.046875,-0.0078125,0.0390625,0.015625,-0.0078125,-0.0078125,-0.0078125,-0.015625,-0.0625,-0.0625,-0.015625,0.0234375,0.078125,0,0.0078125,0.0078125,0.0078125,-0.0078125,-0.046875,0.0234375,-0.0078125,0.0078125,-0.0078125,0.0078125,0.0078125,0,-0.0078125,-0.0078125,0,0.09375,0.015625,-0.0234375,-0.0390625,-0.015625,0.0078125,-0.0546875,-0.078125,-0.046875,-0.0234375,-0.0078125,0.03125,0.1953125,0.0703125,-0.03125,0.0625,0.0078125,0.03125,0.0234375,-0.0390625,-0.0078125,0.1171875,0.0625,0.0078125,-0.015625,-0.0625,-0.046875,-0.0078125,-0.0234375,0,0.015625,-0.015625,0.0078125,0.0078125,-0.0390625,0.015625,-0.015625,-0.046875,-0.0078125,-0.0234375,-0.0546875,-0.015625,0.0546875,0,-0.0234375,0.0546875,0.0078125,0.015625,0.015625,0.015625,-0.0078125,0,-0.03125,-0.015625,-0.03125,-0.0078125,0,0.0234375,0.0703125,0.0078125,-0.015625,0,0.0234375,0.0234375,0.0390625,0.0078125,-0.046875,0.015625,0.015625,-0.0390625,-0.0390625,-0.03125,-0.1015625,-0.1171875,-0.0078125,-0.0390625,-0.0390625,-0.0234375,0.0234375,-0.0078125,-0.0078125,0.0390625,0.0234375,-0.046875,0.0234375,-0.0078125,-0.015625,-0.03125,0.03125,0.0625,-0.015625,0,0.015625,0.0078125,-0.015625,0,0,-0.015625,0.0078125,0.015625,0,-0.0078125,-0.0078125,-0.0546875,0.0078125,0.0234375,0,-0.0234375,-0.015625,-0.0234375,-0.015625,0,0,-0.03125,-0.0078125,-0.0078125,0.046875,0.0546875,-0.0078125,-0.0234375,0,-0.0234375,-0.015625,-0.0546875,-0.078125,0.03125,0.0078125,0,0,0,-0.0234375,-0.015625,-0.0234375,0.046875,0.015625,0,-0.0390625,0.015625,-0.0625,-0.03125,-0.03125,-0.0859375,-0.0625,0.0234375,-0.03125,0,-0.0234375,0.046875,0.015625,-0.0390625,-0.015625,0.046875,-0.015625,-0.015625,-0.0234375,-0.0234375,-0.0625,0.0078125,-0.0078125,-0.0390625,0,0.0546875,-0.0546875,-0.0234375,-0.0078125,-0.0703125,-0.078125,-0.0234375,0.0390625,0.015625,-0.0625,-0.0234375,-0.015625,0,-0.0390625,0.0625,0.0625,-0.0078125,-0.0625,0.0078125,0.0703125,0.0625,0.0234375,-0.078125,-0.0625,0.0234375,-0.0390625,0.0078125,0.0078125,-0.0546875,0.0078125,-0.046875,0.0859375,0.03125,0.03125,0.046875,-0.0078125,-0.046875,-0.015625,-0.046875,-0.0234375,0.0078125,-0.0859375,-0.0234375,-0.0625,0.0234375,0,-0.03125,-0.0234375,-0.0078125,-0.0078125,0,0.0390625,0,-0.015625,-0.0234375,-0.046875,-0.0234375,0.0234375,0.0703125,-0.0078125,-0.046875,0.0390625,0.1171875,0.0390625,-0.0390625,-0.0390625,0,0.03125,-0.0234375,-0.015625,0.109375,-0.0625,0.015625,-0.03125,0.0078125,0,0,-0.0234375,-0.046875,-0.0234375,-0.0625,-0.0859375,0,-0.0078125,0.0078125,0.0078125,0,0.015625,0.0078125,-0.015625,-0.0078125,-0.0078125,0.03125,0.0390625,0.09375,-0.09375,-0.015625,-0.0859375,0.03125,-0.015625,-0.015625,0.015625,0.0078125,0.046875,-0.0703125,-0.046875,-0.03125,-0.0390625,0.078125,-0.03125,-0.015625,0.0078125,-0.09375,-0.03125,0.0859375,-0.0703125,0.0859375,0.140625,0,0.0078125,-0.0078125,0,0.0078125,0,0,0.0078125,0,0.09375,-0.0546875,0.0859375,-0.0234375,0.015625,-0.1328125,-0.03125,0.1328125,-0.09375,-0.0390625,-0.0390625,-0.1015625,-0.03125,0,0.0234375,-0.0390625,-0.03125,0.1328125,0,-0.078125,-0.078125,0.015625,0.125,-0.078125,-0.0859375,-0.0234375,0.0390625,0.03125,-0.0234375,-0.0390625,0.0625,-0.09375,-0.0234375,0.0390625,-0.0078125,-0.015625,0.03125,-0.0546875,-0.0390625,-0.0390625,0.03125,-0.078125,-0.0078125,0.109375,0.1015625,-0.0078125,0.0078125,0.0390625,0,0.078125,0.09375,0.0390625,-0.0234375,-0.0625,0.0234375,0.03125,-0.015625,0.046875,0.0234375,-0.0234375,-0.0078125,0.0546875,-0.015625,0.0078125,-0.015625,0.015625,-0.046875,-0.0703125,-0.03125,-0.0625,0.0390625,-0.0703125,-0.0234375,-0.0546875,0.03125,-0.0078125,0.046875,0.0390625,-0.0703125,-0.0390625,0.0390625,-0.015625,-0.0234375,0.0859375,-0.03125,-0.109375,0.0390625,0.046875,-0.109375,-0.0078125,-0.0078125,0.0078125,0.015625,-0.015625,-0.0234375,0,-0.0078125,-0.0078125,0,-0.03125,-0.0078125,0.015625,0.0703125,-0.0859375,-0.015625,0.03125,-0.0390625,-0.046875,-0.03125,0.0234375,-0.0234375,0.0078125,-0.046875,0.015625,0.0078125,-0.0625,-0.0234375,0.015625,-0.0546875,-0.078125,0.0390625,0.0234375,0.015625,0,-0.015625,-0.015625,-0.015625,-0.0859375,-0.09375,0.0078125,0,0.0859375,0.015625,-0.0078125,0.0078125,0.0234375,-0.015625,0.0234375,0.015625,-0.03125,0.0859375,0,-0.0546875,-0.0546875,-0.015625,0.03125,0.015625,0.0078125,-0.0625,0.03125,0.0234375,0.0078125,-0.0546875,-0.078125,0,0.0546875,0.0703125,0.0078125,0.0546875,0.0234375,-0.03125,-0.0703125,-0.015625,0.0078125,0,-0.0078125,0.0859375,0.015625,0,0.0078125,0.0546875,0,0.0078125,-0.046875,-0.109375,0.015625,-0.0078125,-0.0390625,0.078125,0.078125,0.0546875,-0.015625,-0.0703125,0.09375,-0.0078125,-0.0703125,0.078125,-0.015625,-0.0546875,-0.1015625,-0.078125,0.03125,0.015625,-0.0390625,0.0703125,-0.015625,0.0703125,-0.1875,-0.03125,-0.03125,-0.015625,-0.0546875,-0.0078125,-0.015625,-0.1171875,0.0078125,-0.0234375,0,0,0.0078125,0.0234375,-0.0625,-0.09375,-0.0078125,0,-0.015625,-0.0234375,-0.0546875,-0.078125,0.0703125,-0.015625,-0.0078125,0.0078125,-0.015625,-0.015625,-0.1015625,-0.09375,-0.015625,0.0625,0.015625,-0.0078125,0.1796875,-0.0859375,-0.0234375,-0.015625,0.0703125,0,-0.0390625,0,-0.0859375,-0.015625,-0.0078125,-0.046875,0.0078125,0,-0.0078125,-0.0078125,0.0078125,-0.0078125,0,0.0078125,-0.015625,0.0390625,0.0390625,0.0078125,0,0.0234375,0.0078125,-0.0546875,-0.0625,-0.078125,0,0.03125,-0.015625,0,0.0078125,0.015625,0.0078125,0.0078125,-0.0078125,-0.015625,0.015625,-0.046875,-0.03125,0.0078125,0.03125,0.1015625,0.0234375,-0.015625,-0.0078125,-0.0078125,0,0,0.0078125,0.0078125,-0.0078125,-0.015625,-0.0078125,-0.015625,0,-0.0078125,-0.0390625,-0.0234375,-0.03125,-0.0234375,0.046875,-0.0390625,-0.0546875,-0.078125,0.0625,0.015625,-0.0546875,-0.078125,0.1015625,-0.09375,-0.0390625,0.015625,0.0390625,0.078125,0,-0.078125,0.03125,-0.03125,0.0234375,0.03125,0.0234375,0.0078125,0.0078125,0.03125,0.046875,-0.015625,-0.0078125,-0.046875,-0.046875,-0.0078125,0.0234375,0.0390625,-0.046875,-0.0234375,-0.0546875,0.0234375,0.125,-0.0078125,-0.0078125,0.0078125,0.0078125,0.015625,0.0546875,-0.0390625,-0.0390625,-0.03125,0,0.015625,-0.03125,0.0234375,0.0078125,-0.0234375,0,0.0234375,0.0078125,0.015625,0,-0.0234375,0.0078125,-0.0234375,-0.03125,0.09375,-0.03125,0.0390625,0.015625,0.0078125,-0.046875,-0.03125,-0.0546875,0.09375,0.0390625,-0.0234375,-0.0625,0.0078125,0.03125,-0.0703125,0.0078125,-0.0390625,0.03125,-0.1015625,-0.0546875,0.0703125,0,0.015625,0.0078125,0,0.0078125,-0.015625,-0.015625,-0.0078125,-0.0078125,0,-0.0078125,0.046875,-0.0078125,-0.015625,-0.0390625,-0.03125,-0.0078125,-0.0234375,0.0078125,-0.0390625,-0.0625,-0.046875,-0.015625,0.1171875,-0.0078125,0.0078125,-0.0078125,-0.0703125,-0.03125,-0.046875,0.015625,-0.046875,-0.0234375,0.0078125,-0.046875,0,-0.0078125,-0.03125,0.0078125,-0.0390625,-0.0390625,0.0234375,0.015625,-0.03125,0.046875,0.015625,0.046875,-0.015625,-0.046875,0.0390625,0.0234375,-0.03125,-0.0078125,-0.03125,-0.078125,0.015625,-0.0234375,-0.1015625,0.015625,-0.03125,0,0,-0.046875,-0.0703125,-0.0390625,-0.0625,-0.015625,-0.03125,-0.046875,0.1015625,-0.0234375,-0.015625,-0.046875,-0.015625,0,0.0078125,-0.0390625,-0.015625,-0.0703125,0.03125,0.0234375,-0.0703125,-0.0078125,-0.03125,-0.0625,0.0234375,0.046875,-0.0234375,0.0390625,-0.015625,-0.0078125,0.015625,-0.03125,0.0390625,-0.015625,-0.0234375,0.0625,-0.0390625,-0.0546875,-0.0234375,-0.0078125,0,-0.0546875,0,0.046875,0.078125,0.03125,0.0078125,0.0546875,-0.0546875,-0.09375,-0.0390625,-0.015625,-0.015625,0.109375,0.0078125,0,-0.0390625,-0.015625,0,0.0390625,0.0078125,-0.03125,-0.046875,0.015625,0.015625,-0.046875,-0.03125,-0.0234375,-0.046875,0.03125,-0.0390625,-0.03125,-0.0078125,0.015625,-0.015625,-0.03125,-0.015625,0.078125,0.0078125,0.015625,-0.046875,0,-0.0234375,-0.0078125,-0.0625,0.0859375,0.03125,-0.03125,-0.03125,-0.0234375,0.0234375,-0.0546875,-0.09375,0,-0.0078125,-0.0078125,-0.0078125,0.0078125,-0.015625,-0.015625,0,0.0078125,0,0.046875,0.109375,-0.0078125,-0.0546875,0.0234375,-0.046875,0.0234375,0.03125,-0.03125,-0.0234375,0,-0.0546875,-0.0703125,0.0546875,-0.015625,0.0078125,0.0859375,0.0234375,-0.0859375,0.0078125,0.015625,-0.078125,-0.015625,-0.0390625,0.171875,-0.0390625,0.0078125,-0.0078125,-0.015625,0.0078125,0,-0.0078125,0.0078125,0,0.0078125,-0.046875,-0.046875,-0.0859375,-0.1015625,-0.046875,0.03125,0.03125,-0.0078125,0.03125,0.09375,-0.0234375,-0.03125,-0.0390625,-0.0078125,-0.0078125,-0.0234375,0,-0.0546875,0,-0.0078125,0,-0.0078125,0.015625,0.0859375,-0.0078125,0.0546875,-0.1015625,-0.046875,-0.03125,0.078125,0.03125,-0.015625,-0.0234375,0,-0.0234375,-0.015625,0.015625,-0.015625,-0.0625,-0.0546875,-0.015625,0.078125,-0.0703125,-0.0546875,-0.0390625,-0.0078125,-0.03125,-0.015625,-0.0078125,0,0.0078125,-0.015625,-0.03125,-0.0546875,0.015625,-0.0078125,-0.015625,-0.0234375,0.0078125,0.0078125,0.046875,0.03125,0.0078125,0.0078125,-0.015625,-0.0625,-0.0078125,0.0234375,0.046875,-0.046875,0.0078125,-0.015625,-0.0078125,0.0625,0.046875,-0.015625,-0.0390625,0.0234375,0.015625,-0.15625,-0.046875,-0.0234375,-0.0234375,0.0703125,0.0390625,-0.015625,-0.03125,0.015625,0.0234375,0.03125,0,0.0078125,0,-0.015625,-0.015625,0,-0.0078125,0.015625,0.0078125,0,-0.0546875,-0.0078125,0.0234375,-0.0546875,-0.0390625,-0.0390625,0.046875,-0.0078125,0.0078125,-0.0078125,-0.0390625,0.03125,0.0625,0.0625,-0.015625,-0.046875,0.0546875,0.03125,0,0.03125,-0.03125,0.015625,0.0234375,0.0546875,-0.0234375,-0.0234375,0.0078125,-0.03125,0,0.0390625,-0.015625,0.046875,-0.1015625,-0.0625,0.015625,-0.046875,-0.03125,0.0234375,-0.0078125,0.015625,0.046875,-0.0234375,0.0078125,0.0234375,-0.03125,0.0078125,-0.0234375,-0.0625,0,-0.015625,-0.0234375,0.015625,0,0.046875,-0.0703125,-0.0703125,-0.0390625,0.0703125,0.0078125,0,-0.015625,0.0234375,-0.0078125,-0.0234375,-0.015625,0.03125,-0.078125,-0.015625,-0.0078125,0.0234375,-0.0078125,0.0234375,0.0390625,0.0546875,-0.046875,-0.0546875,-0.0078125,-0.015625,0.046875,-0.0546875,0.0546875,0.0390625,-0.046875,0.0078125,-0.0546875,0.046875,0,0.0390625,-0.0234375,-0.0078125,-0.0234375,0,0.0546875,0.109375,0.0078125,-0.0078125,-0.046875,-0.0078125,0,-0.0390625,0.0234375,-0.0546875,-0.0234375,0.0078125,-0.046875,0.015625,-0.046875,0.03125,-0.0078125,-0.03125,-0.0859375,-0.0703125,0.015625,-0.0234375,-0.015625,0.0859375,0.0625,0.0078125,-0.0703125,0,-0.046875,0.0078125,0.0390625,-0.0234375,0.03125,0.0234375,-0.0234375,0.0234375,0.0390625,0,0,0,0.0234375,0.0859375,-0.03125,-0.03125,0,0.125,-0.0390625,0,-0.0546875,-0.0625,0.015625,0,-0.0078125,-0.015625,-0.0078125,0.0234375,0.0078125,0.0078125,0.0078125,0.0078125,0.0390625,-0.0234375,0.015625,0,0.03125,0.0234375,-0.015625,-0.0625,0.03125,-0.0234375,-0.0625,-0.03125,0.1171875,-0.0234375,-0.015625,0.0546875,-0.0078125,0.0859375,-0.03125,0.078125,0.0234375,0.0234375,-0.03125,-0.015625,0.078125,0.0546875,0.0625,0,-0.0078125,0.0078125,-0.015625,-0.0078125,-0.0078125,-0.0078125,0,0,0.0390625,0.0546875,-0.0078125,0.1171875,-0.0078125,-0.0546875,-0.109375,0.0703125,0.046875,0.0078125,-0.046875,-0.0078125,-0.0078125,0.015625,-0.0390625,-0.0390625,-0.015625,0.0625,0.078125,0.0078125,-0.03125,0,-0.0078125,-0.078125,-0.0546875,-0.046875,0.078125,0.0078125,-0.046875,0.0078125,0.0390625,0.015625,0.0078125,0.0078125,-0.078125,-0.03125,0,-0.0078125,-0.015625,-0.046875,-0.0546875,-0.0078125,0.0859375,-0.03125,-0.015625,0.0234375,0.015625,-0.0078125,-0.0546875,0,-0.0078125,-0.015625,-0.0234375,-0.03125,0.03125,-0.015625,-0.015625,0.03125,-0.015625,-0.015625,-0.0390625,0.015625,-0.015625,-0.0234375,0,0.0234375,-0.0546875,0.03125,-0.015625,0.046875,-0.0234375,-0.015625,-0.0234375,0.0078125,-0.015625,0.0546875,-0.046875,-0.0859375,0.0390625,-0.0625,-0.03125,-0.0234375,0.0234375,-0.0625,-0.078125,0.015625,0,0.0859375,-0.0390625,0.0078125,0.0078125,0.0078125,0,0,-0.0078125,-0.0234375,0.0078125,-0.0078125,0.0078125,-0.0234375,0.0390625,0.0078125,0,-0.015625,0.0234375,0.0078125,0.0078125,0.0078125,-0.03125,-0.03125,-0.0078125,0.125,-0.078125,0.0390625,-0.0390625,-0.0234375,-0.015625,0.0078125,-0.03125,0.0078125,-0.03125,0.0234375,-0.0234375,-0.015625,0.0390625,-0.0546875,0.03125,-0.03125,-0.03125,-0.078125,-0.0703125,-0.015625,0.078125,0.03125,-0.078125,-0.03125,-0.015625,-0.015625,-0.0625,-0.078125,0.03125,0.0703125,0.0625,0,-0.015625,0.015625,0,0.0703125,-0.0390625,-0.015625,-0.0703125,-0.046875,-0.046875,-0.0625,-0.09375,0.015625,-0.03125,-0.0625,0.03125,0.1171875,0.0390625,-0.0625,0.0546875,0.0078125,-0.0078125,0.015625,0.0078125,-0.0390625,0,0.0078125,0.0078125,-0.046875,-0.0625,-0.03125,-0.03125,-0.0234375,0.046875,0,-0.0703125,0.046875,0.015625,-0.0390625,-0.015625,0,0.0234375,-0.03125,-0.0859375,0.046875,-0.03125,0,0.0625,0.0234375,0.015625,-0.03125,-0.078125,0.125,-0.0703125,-0.0078125,-0.0859375,0.0078125,-0.0078125,0.046875,0.046875,-0.09375,0.0625,0.125,-0.0390625,-0.046875,-0.0234375,-0.03125,0,-0.03125,-0.0546875,0.0390625,-0.078125,-0.015625,-0.015625,-0.0234375,-0.03125,0.0859375,-0.015625,-0.046875,-0.0859375,-0.0546875,0.0625,-0.0625,-0.0234375,-0.015625,0.0234375,-0.03125,-0.015625,0.046875,-0.0234375,-0.0546875,-0.0390625,0.0625,-0.078125,-0.0546875,0.0234375,-0.0078125,-0.0390625,0.0078125,-0.046875,-0.0078125,0,0,0.0078125,0,0,0,-0.0078125,-0.015625,-0.0078125,-0.015625,0.0078125,0.0078125,-0.0859375,0.0546875,-0.0390625,-0.078125,0.0625,-0.03125,-0.078125,0.078125,0.03125,0,-0.1171875,-0.0546875,-0.03125,0.0859375,-0.015625,0.015625,-0.0078125,-0.03125,-0.0859375,0.0390625,-0.0234375,-0.09375,0.0390625,-0.015625,0.0078125,0,-0.0078125,0,0.0078125,0.0078125,0,-0.015625,0.0546875,0,0.046875,-0.03125,0.0546875,-0.09375,-0.03125,-0.0234375,-0.0625,0.0625,-0.015625,-0.1015625,0.03125,-0.078125,0.0703125,-0.0703125,-0.015625,0,-0.0234375,-0.015625,-0.0703125,-0.0546875,0.0390625,0.046875,-0.0234375,-0.0546875,0.109375,-0.03125,0.0234375,-0.03125,0,-0.046875,-0.0078125,0.0078125,0.046875,-0.0234375,-0.0234375,0.046875,0.046875,-0.0390625,0.046875,-0.015625,-0.046875,0.03125,0.015625,-0.015625,-0.0078125,-0.0546875,0.015625,0.0703125,0.0234375,0.0078125,-0.0234375,0,0.015625,-0.0078125,-0.0078125,0.015625,0.0546875,0.015625,0.0078125,-0.015625,-0.046875,0.015625,-0.0390625,0.0859375,-0.03125,-0.078125,0.046875,0.046875,-0.046875,0,-0.0078125,0.015625,-0.0625,-0.0703125,0.03125,0.0234375,0.0390625,-0.015625,0.015625,-0.0390625,0.1015625,0.0234375,-0.0234375,-0.0703125,0.1015625,0.0625,-0.03125,-0.0078125,-0.015625,-0.03125,-0.015625,-0.015625,0,0.0234375,-0.0078125,0.015625,0.0390625,0,-0.0234375,-0.0390625,0.0078125,-0.0078125,-0.015625,-0.0078125,0.03125,0.03125,-0.078125,-0.015625,0.0078125,0.015625,-0.046875,-0.015625,-0.03125,-0.0234375,-0.015625,0.0546875,0.0234375,-0.0546875,0.0078125,-0.0546875,0.0625,0.0234375,0.03125,0.0234375,-0.0078125,0.0390625,-0.0390625,0.0078125,-0.046875,-0.0078125,0.03125,0.0859375,-0.0390625,-0.0078125,-0.0078125,-0.0703125,-0.015625,0,-0.0625,-0.0390625,0.0234375,0.0234375,-0.0390625,-0.0625,-0.09375,-0.0390625,-0.0546875,0.0234375,-0.0234375,0.0390625,0.078125,0.0390625,-0.0703125,0.046875,0.0234375,-0.09375,0.09375,-0.0234375,0.0078125,0.140625,-0.03125,0.03125,-0.0703125,0,-0.0703125,0.0234375,0,0,0.015625,-0.0078125,0,0.03125,-0.0625,-0.0390625,0.1171875,0,-0.0078125,0.0078125,0.0703125,-0.0546875,0.0078125,0.0390625,0.0234375,0.0078125,-0.0625,-0.015625,0.1484375,-0.078125,0.0234375,0.1328125,-0.0390625,-0.1640625,0.109375,0.1171875,0.03125,-0.0703125,-0.0390625,0.0234375,0.0234375,-0.015625,0.0234375,-0.046875,-0.0546875,-0.0078125,-0.0390625,-0.015625,-0.109375,0.09375,0.0703125,-0.0859375,-0.03125,-0.0546875,-0.0390625,0.03125,-0.015625,-0.0546875,-0.0625,0.0546875,-0.09375,0.0625,-0.046875,-0.0546875,0.0234375,-0.0078125,0.046875,0,-0.03125,0.03125,-0.03125,-0.1015625,-0.0390625,-0.0546875,0.0078125,0.0078125,-0.0234375,-0.015625,0.03125,0,-0.0390625,-0.0078125,0.015625,0.0078125,0.0078125,-0.0078125,-0.0078125,-0.015625,0,0,0.0078125,-0.0078125,0.0234375,-0.0234375,-0.0078125,0.046875,0.015625,0.015625,-0.0078125,-0.0234375,-0.0390625,0,0.03125,-0.03125,0.03125,-0.03125,0.03125,0.0234375,-0.03125,-0.0234375,0.0390625,0.03125,0.03125,0.0390625,-0.0078125,-0.0078125,-0.0234375,-0.0078125,-0.0078125,0,0,0.0078125,-0.015625,0,-0.0078125,0,0.0078125,-0.0078125,0.0234375,0.0234375,0.015625,0.0390625,-0.0390625,-0.0234375,-0.0390625,-0.046875,0.0625,-0.015625,0,0.0234375,0.015625,-0.0078125,-0.015625,0.0390625,-0.0234375,-0.015625,0.0234375,-0.0078125,-0.015625,0.015625,-0.0625,0.078125,-0.0390625,-0.046875,0.015625,-0.03125,-0.03125,-0.0234375,-0.015625,0.0078125,0.0625,0,-0.0390625,0.0078125,-0.0078125,0,0,-0.03125,0.0078125,0.078125,-0.03125,-0.0078125,-0.0078125,-0.0390625,0.0078125,0.0078125,-0.015625,0,-0.0234375,-0.0078125,0.015625,-0.0234375,-0.0234375,0.0078125,0,0.0078125,0.0078125,-0.0234375,0,0,0.0078125,0,0.0078125,-0.0234375,-0.015625,0.015625,-0.015625,-0.0234375,-0.015625,0,0.046875,0.0390625,-0.015625,-0.0234375,0.0078125,0.0234375,-0.015625,-0.0625,0.0234375,0.03125,-0.03125,-0.0078125,0.015625,0.0078125,0.015625,0.0078125,-0.015625,0.015625,0.0234375,0.0234375,-0.0078125,0,0,-0.0078125,0,-0.0078125,0.0078125,-0.03125,-0.015625,-0.0234375,0,-0.0390625,-0.03125,0.015625,0,-0.0078125,-0.0078125,-0.0390625,0.0078125,0.015625,-0.015625,-0.015625,0,-0.0390625,0.0078125,-0.03125,-0.078125,0.0234375,0.0703125,0,-0.0078125,0.0234375,-0.0234375,0.015625,0.0234375,-0.0078125,0.0078125,0.0703125,0.046875,-0.0234375,-0.0078125,-0.0078125,-0.046875,0.015625,0.03125,0.0078125,-0.0546875,-0.078125,-0.03125,0.0078125,-0.0234375,0.03125,0.0234375,-0.0078125,0,0.03125,0.015625,-0.0390625,-0.03125,-0.0234375,-0.046875,-0.0390625,-0.046875,-0.0234375,0.0625,0.03125,0,0,0.015625,-0.0234375,-0.0390625,-0.015625,0,0.046875,-0.0234375,-0.015625,0.0078125,-0.03125,-0.015625,0.0234375,0.0390625,-0.015625,-0.015625,0,-0.078125,-0.0234375,-0.0078125,-0.03125,-0.03125,0.015625,0,0.0390625,0.03125,-0.0078125,-0.0234375,-0.0078125,-0.0234375,-0.0546875,0.015625,-0.078125,-0.03125,0.015625,0.0390625,-0.0390625,-0.0546875,-0.0234375,0,-0.046875,0,0.0234375,-0.0234375,0.0234375,0,0.015625,0.0546875,0.0234375,-0.0390625,0,0.046875,0.046875,0.0078125,0,-0.0390625,-0.015625,-0.0390625,-0.046875,0.015625,0.0625,0.0703125,-0.0078125,-0.0078125,0.015625,0.03125,-0.0234375,-0.0234375,0.0078125,0.0390625,0.046875,-0.0234375,0.0234375,-0.0078125,-0.03125,0.0234375,0.0078125,-0.015625,0.015625,-0.0546875,-0.0390625,-0.0390625,-0.0546875,-0.046875,0,-0.015625,0,0.0078125,0,0.015625,0.0078125,0,-0.0078125,0.0078125,-0.0234375,-0.015625,0.0390625,0.0625,-0.0546875,0.015625,-0.0078125,0.0234375,-0.015625,0.0546875,-0.015625,0.0234375,-0.015625,0,0.03125,-0.078125,0.0390625,-0.0078125,0.0390625,-0.0390625,-0.03125,0.015625,0.078125,0,-0.0390625,0.015625,0,-0.0078125,-0.0078125,0,-0.0078125,0.0078125,-0.0078125,0.0078125,0,-0.0390625,-0.0625,-0.0390625,0.015625,0.0625,0.015625,0.0390625,-0.046875,0.078125,-0.078125,0,0.0078125,0.078125,0.078125,-0.03125,0.0625,0.0078125,0.0234375,-0.03125,0.0390625,-0.078125,0.015625,0.03125,0.015625,0.03125,-0.0625,-0.0390625,0.0078125,-0.015625,0.0078125,0.0078125,0.0390625,0,0.0390625,0.0234375,0.0625,-0.0078125,0,-0.03125,-0.078125,-0.0546875,-0.109375,0.046875,0.015625,0.0703125,0.0234375,0.078125,-0.0078125,-0.0234375,-0.0234375,0.0078125,-0.0234375,0.0234375,-0.0234375,-0.0234375,-0.0390625,0.03125,0.03125,0.015625,0.0078125,-0.0234375,-0.015625,0.015625,0.015625,0.03125,0.0703125,-0.03125,0.015625,0.015625,-0.0546875,-0.0234375,-0.0390625,0.0390625,-0.046875,0.0078125,-0.0078125,-0.015625,-0.0078125,-0.0625,-0.0859375,-0.03125,0.046875,-0.046875,-0.046875,0.0546875,-0.03125,0.0390625,0.0234375,-0.046875,0.0546875,0.0078125,0,-0.015625,0.015625,-0.0078125,0,0.0078125,-0.0234375,-0.015625,-0.015625,0.0859375,0.03125,-0.015625,-0.03125,-0.03125,0.03125,0.0234375,-0.03125,-0.046875,-0.0390625,0.03125,-0.0078125,0,-0.015625,0.03125,0.0234375,-0.0546875,-0.0078125,-0.0234375,0,-0.0546875,0.0546875,-0.0078125,0.0234375,0.0546875,-0.0625,0.015625,0.0078125,-0.0703125,-0.046875,0.0546875,0.0078125,0.015625,-0.0703125,0.03125,0.0546875,0.015625,-0.0078125,0.078125,0.0078125,-0.0703125,0.0078125,0,-0.0625,0.015625,0,0.046875,0.078125,-0.0078125,0.03125,0.03125,-0.0390625,-0.0078125,-0.0390625,-0.1015625,0.1171875,-0.0390625,-0.0859375,0.0703125,0.046875,-0.046875,-0.015625,0.0625,0.09375,0.015625,0.0078125,-0.015625,-0.046875,-0.03125,-0.03125,0.0234375,0.03125,0.03125,0.0078125,0.0234375,-0.0234375,-0.0546875,-0.03125,0.09375,-0.015625,-0.015625,-0.0078125,0,0.0390625,0.0234375,-0.0078125,-0.03125,-0.03125,0,-0.0703125,0.0625,0,-0.015625,-0.0390625,-0.03125,-0.0390625,-0.0703125,0.0390625,0.0625,-0.03125,-0.0625,-0.015625,-0.046875,-0.046875,0.015625,0.015625,0.0078125,0,-0.0390625,-0.0078125,-0.0390625,-0.015625,-0.03125,0.0234375,0.046875,0,0.0078125,-0.015625,0.0703125,0.0390625,0,0.0625,-0.03125,0.0078125,-0.03125,-0.046875,0.015625,0.0390625,-0.0859375,-0.0078125,-0.0546875,0.0390625,0.046875,-0.0390625,-0.0078125,-0.015625,-0.03125,0.0390625,0.0234375,0.0078125,0,0.03125,0.0703125,0,-0.015625,-0.015625,0,0,0.015625,0,-0.015625,0,0.0390625,-0.03125,-0.078125,-0.0234375,-0.015625,-0.0234375,-0.0390625,0.1015625,0.0859375,0.0078125,-0.0390625,0.03125,-0.015625,0.03125,-0.0234375,-0.0078125,-0.0390625,0.0234375,0.03125,-0.0078125,-0.0625,-0.078125,0.015625,0.0234375,-0.046875,-0.0390625,0.0390625,0,0.0078125,0.0078125,-0.0078125,-0.0078125,0,0.0078125,0,-0.015625,0.046875,-0.0625,-0.0625,-0.03125,-0.046875,0.0625,-0.046875,-0.0625,0.0703125,-0.1015625,0.0546875,-0.0546875,-0.046875,0.015625,0.0390625,0.0390625,-0.0078125,0.0078125,-0.0390625,-0.046875,-0.0234375,0.0859375,0.0390625,-0.015625,-0.0234375,-0.015625,-0.078125,0.0078125,0.0078125,-0.015625,-0.03125,-0.015625,-0.046875,-0.046875,0.0390625,0.0390625,0.109375,0,0.0625,0.0078125,-0.0703125,-0.0703125,-0.0390625,-0.015625,0.0234375,-0.0390625,0.0390625,-0.0078125,-0.0078125,-0.0390625,-0.0390625,0,-0.0625,0.0078125,-0.0078125,-0.03125,-0.0078125,-0.0078125,0.0078125,0.046875,0,0,0.0234375,-0.015625,-0.0078125,0.0234375,-0.015625,-0.1328125,0.125,-0.015625,-0.03125,-0.0078125,0.1015625,0.0234375,-0.078125,-0.015625,-0.1015625,-0.03125,0.0703125,-0.03125,-0.015625,0.0859375,0.0390625,-0.0625,0,-0.0390625,0.0234375,0,-0.0546875,0.0859375,0,-0.0078125,-0.015625,0.0078125,0,0.015625,0.015625,0,0.0234375,0.0078125,0.0390625,-0.0546875,-0.0078125,0.015625,0.0234375,0.0078125,0.0078125,-0.0078125,-0.078125,0.0625,0.0703125,-0.0625,-0.078125,-0.015625,-0.0390625,0.0234375,0.0546875,-0.046875,0.046875,-0.0546875,-0.0625,-0.0703125,-0.015625,-0.0390625,0.0078125,0.1328125,-0.0234375,0.015625,-0.1328125,-0.0078125,-0.1484375,-0.0703125,0.0546875,0.0390625,0.0859375,0.0703125,0.0625,-0.0390625,0.0234375,-0.0703125,-0.0625,-0.015625,-0.0078125,0.0859375,0.03125,-0.0703125,-0.0390625,0.0625,0.0390625,0.0546875,0.0078125,0.0546875,-0.0078125,-0.0546875,-0.0390625,0.15625,-0.1015625,-0.125,0.046875,0.046875,-0.015625,0.0234375,-0.015625,0.0390625,-0.09375,-0.0078125,0.0078125,-0.1328125,0.015625,0.046875,-0.0234375,-0.0078125,0.03125,0.0234375,-0.03125,-0.078125,0.0625,0.0546875,-0.0859375,0,-0.0390625,-0.0859375,-0.0625,-0.0390625,-0.03125,0.0859375,-0.015625,-0.078125,0.140625,-0.046875,0,0.0546875,-0.109375,-0.1875,-0.0234375,0.015625,-0.0390625,-0.0625,0.0234375,0.1015625,0,-0.0546875,0.0078125,0.03125,-0.03125,0.0859375,0.0078125,0.046875,-0.0625,0.1171875,-0.0234375,-0.109375,0.03125,-0.0625,-0.0234375,-0.0625,-0.0390625,-0.09375,0.0234375,-0.015625,0.0234375,0.0625,-0.0078125,-0.015625,0,0.015625,-0.0234375,0.0625,0,-0.078125,0,-0.0859375,0.078125,0.03125,0.0390625,-0.0390625,-0.0859375,-0.03125,0.03125,0.0703125,0.0234375,-0.03125,-0.0234375,0.015625,0.0078125,0.0078125,0,-0.0078125,-0.0078125,0.0078125,0,-0.0078125,0.03125,-0.03125,-0.078125,-0.0546875,-0.078125,0.0078125,0.015625,-0.015625,0.03125,0,-0.09375,-0.046875,0.03125,-0.03125,-0.015625,0.0234375,-0.046875,0,0,-0.0625,0.0546875,0.140625,-0.09375,0.03125,0.0390625,0,-0.078125,-0.0234375,0,0,0.0078125,0.015625,-0.015625,-0.0078125,0.0078125,0,-0.0234375,-0.0390625,0,-0.0078125,0.0390625,-0.078125,0.015625,0.015625,0.03125,-0.0703125,0.046875,-0.046875,-0.0859375,-0.0546875,0.078125,-0.0546875,0.0078125,0.03125,0.015625,0.046875,0.0234375,0.03125,0.0078125,0,0,-0.0703125,-0.0390625,0.046875,0,-0.03125,0.0078125,0.0234375,-0.015625,-0.0234375,-0.0078125,-0.015625,0.0234375,0.046875,0.0234375,0.0234375,0.0703125,0.0078125,-0.0234375,0.0390625,0.0546875,0.0390625,-0.015625,0.0078125,0.0078125,-0.046875,-0.0234375,0,0.015625,0,-0.015625,-0.015625,-0.0234375,-0.015625,0,0.0078125,-0.046875,0.015625,0,0,-0.0390625,-0.0390625,0.0703125,0.015625,0,-0.0390625,-0.046875,0.015625,-0.015625,-0.0390625,-0.0390625,0.046875,0.15625,-0.015625,-0.015625,-0.015625,0.0625,-0.078125,0.078125,-0.015625,-0.0859375,0.046875,-0.03125,0.0625,0.0234375,0.0234375,-0.015625,-0.0078125,-0.0078125,0,0.0078125,0,-0.015625,0.015625,-0.0078125,-0.015625,-0.0234375,0,-0.015625,-0.03125,0.0546875,0,0,0.0390625,-0.0390625,-0.0625,-0.0546875,0.0078125,-0.03125,0.0703125,-0.0625,-0.0234375,-0.03125,-0.0390625,-0.0078125,-0.0078125,0.0703125,0.0078125,0.0078125,0.0546875,0.09375,-0.0234375,-0.046875,-0.0859375,-0.0703125,0.0234375,0.015625,0.03125,-0.0859375,-0.0078125,0.03125,-0.0078125,-0.0625,-0.0078125,-0.0390625,0,0.0078125,-0.03125,-0.0390625,-0.0390625,0.0234375,-0.03125,-0.0546875,0.015625,0,-0.03125,-0.0390625,0.046875,-0.015625,0.078125,0.0234375,-0.0859375,0.046875,-0.0546875,-0.0234375,-0.0390625,-0.0234375,-0.0078125,0.015625,0.0546875,0.078125,-0.015625,0.03125,-0.0234375,-0.09375,0,0,-0.0078125,-0.046875,-0.0078125,0.03125,-0.0703125,0.1015625,-0.0390625,-0.0859375,-0.046875,-0.015625,-0.0703125,0,0.078125,0.0234375,0.03125,0.0625,0.015625,-0.03125,0.0703125,-0.0390625,-0.078125,-0.0078125,0.0234375,-0.0234375,-0.0546875,-0.09375,0.0078125,0.09375,0,-0.03125,-0.0234375,0,-0.03125,-0.015625,-0.03125,0.03125,-0.0078125,0.0234375,-0.0546875,-0.015625,-0.078125,0.0234375,-0.015625,-0.0390625,0.015625,0.0625,-0.03125,-0.03125,-0.078125,-0.09375,-0.0390625,0.0078125,0.03125,0,0.03125,-0.0078125,-0.03125,-0.046875,0.0078125,-0.015625,0.0390625,-0.03125,0.0078125,0.03125,0.0625,-0.015625,0.0625,0.015625,0.046875,0.0390625,-0.0234375,0,0,0.015625,0,-0.015625,-0.0234375,-0.0078125,0.0078125,-0.015625,-0.015625,0.0078125,-0.1171875,-0.0546875,0.046875,-0.0703125,-0.03125,-0.0703125,0.0390625,0.046875,-0.046875,-0.03125,-0.0546875,-0.0390625,-0.125,0.0703125,0.046875,0.0859375,0.1640625,-0.0546875,-0.0703125,-0.015625,0.0390625,-0.078125,0.1015625,-0.0390625,-0.0703125,-0.0703125,0.0078125,0,0,0.0078125,0,-0.0078125,-0.0078125,0.0078125,0,0.0234375,-0.046875,0.0625,0.15625,0.1015625,-0.078125,-0.1171875,0.015625,0.0546875,-0.0234375,-0.0703125,-0.0078125,-0.015625,-0.0546875,0.0546875,0.0078125,-0.015625,0,-0.0234375,-0.0390625,0.0234375,-0.046875,-0.0703125,-0.0078125,-0.046875,0.0234375,0.140625,-0.03125,-0.09375,-0.046875,-0.046875,0.03125,0.03125,0.0234375,0.0078125,0.0078125,0.046875,0.046875,0.046875,0.0390625,0.0234375,0.140625,0.03125,0,0.0625,0.0234375,0.046875,0.046875,-0.015625,-0.0078125,0.0390625,0.0703125,-0.046875,-0.0390625,-0.015625,-0.0078125,0.0078125,0.0625,-0.015625,-0.03125,0.0078125,0.03125,-0.0078125,0.0390625,0.015625,0,0.0546875,0.0546875,-0.0625,0.0078125,-0.03125,-0.0859375,-0.015625,-0.015625,0.0234375,-0.03125,-0.09375,-0.0078125,-0.0390625,0.0703125,0.078125,0.015625,0.03125,-0.015625,0.0546875,-0.03125,-0.09375,-0.0625,-0.0234375,-0.125,0.015625,0.0234375,0,0.015625,0.0234375,0.0234375,-0.03125,0,-0.0078125,0.015625,0.046875,0,0.0078125,-0.0625,-0.0859375,0.0234375,0.03125,0.0078125,-0.0234375,-0.0859375,-0.0234375,-0.09375,-0.109375,0.1015625,0.0625,-0.0234375,0.09375,-0.03125,-0.0390625,0.0390625,0.0390625,0.0625,-0.0078125,-0.03125,-0.0625,0,0.03125,0.0234375,0.046875,-0.015625,-0.0703125,-0.0078125,-0.0390625,-0.015625,-0.0390625,-0.0234375,-0.0546875,-0.109375,0.0703125,-0.0078125,0.046875,-0.015625,-0.09375,0.0546875,-0.0390625,-0.046875,0.0546875,0.0625,-0.0390625,0.03125,-0.0078125,0.03125,-0.0078125,-0.078125,0.046875,0.1875,0,-0.1796875,-0.0234375,0.0234375,-0.03125,-0.0703125,-0.0234375,0.03125,0.015625,-0.0390625,0.015625,0.0546875,0.046875,-0.03125,0,0.015625,-0.0390625,0,0.0078125,-0.046875,-0.03125,-0.0078125,-0.046875,-0.0859375,0.0078125,-0.09375,-0.0625,-0.03125,-0.0078125,0.03125,0.0078125,0.046875,-0.0078125,-0.078125,-0.1015625,0.0234375,-0.0390625,0.0390625,-0.0546875,-0.0234375,-0.078125,-0.03125,-0.1328125,-0.1015625,0.0546875,-0.0546875,-0.0859375,-0.015625,-0.015625,0.09375,0.0625,0,-0.015625,-0.0390625,0.03125,-0.0390625,0.015625,0.0078125,0.046875,0.1328125,0.015625,-0.0234375,-0.0390625,0.015625,-0.1640625,0.0234375,0.0625,0.0234375,0.046875,-0.046875,-0.0078125,0.0078125,0.03125,-0.109375,-0.0390625,0.0078125,-0.0390625,-0.015625,-0.0546875,-0.1015625,-0.0390625,-0.0625,-0.0703125,-0.0703125,0,-0.0078125,-0.0078125,-0.0078125,0.0078125,0.0078125,0,0,0.0078125,-0.0078125,-0.0234375,0.015625,-0.0078125,-0.015625,0,0,-0.0546875,0,-0.0078125,0.03125,-0.0234375,-0.0234375,0.0546875,-0.015625,0.015625,-0.109375,-0.0078125,-0.03125,0.0546875,-0.0546875,-0.0078125,0.1015625,-0.0234375,0.015625,0.03125,-0.046875,0.0703125,-0.0546875,-0.0625,0,-0.015625,0.0078125,0.015625,0,0.015625,-0.015625,-0.0078125,0.015625,-0.0078125,0.03125,0.0078125,-0.0390625,0,-0.0859375,0.078125,0,0.0546875,0.03125,-0.1328125,-0.0546875,0.03125,-0.0546875,0.0234375,0,-0.0078125,0.0078125,-0.03125,-0.03125,-0.0625,0.0078125,0.125,-0.0390625,-0.0703125,0.1328125,0,-0.0078125,-0.046875,0,-0.0234375,0.0078125,0.03125,0.03125,0.046875,0.0390625,-0.0078125,-0.015625,0.0625,-0.0234375,0.046875,-0.0625,-0.03125,0.015625,-0.015625,-0.1015625,-0.0234375,0.0234375,0.0703125,-0.078125,0.0390625,0.03125,0.0078125,0.09375,0.03125,-0.0234375,0.015625,0.046875,-0.03125,-0.015625,-0.0078125,-0.03125,-0.03125,0.09375,0.0390625,0,-0.015625,-0.0078125,-0.0078125,-0.03125,-0.0078125,0.046875,0.0546875,-0.0625,0.015625,-0.015625,0.03125,0.0234375,0.0234375,-0.046875,0.046875,-0.09375,0.140625,-0.015625,-0.0546875,0.046875,0.1015625,0.0390625,-0.1015625,0.0078125,0.0078125,-0.0078125,0.0078125,0.015625,-0.0078125,0.015625,0,-0.03125,-0.0078125,0.015625,-0.1015625,0.046875,-0.015625,-0.0703125,-0.0546875,-0.03125,-0.0078125,-0.0078125,-0.0078125,-0.046875,-0.0078125,0.0546875,-0.0703125,-0.015625,-0.0078125,-0.046875,-0.0390625,-0.109375,0.0078125,-0.0625,-0.03125,0.0625,0.0234375,0.0234375,-0.0703125,0.0390625,0.015625,0.015625,0.0390625,0,-0.046875,0.0390625,-0.015625,-0.078125,-0.03125,0.03125,-0.015625,0.046875,0,-0.0625,0.015625,-0.0859375,-0.125,0.109375,-0.015625,0.015625,-0.015625,0.03125,-0.046875,-0.0390625,0.078125,0.0703125,-0.0234375,-0.03125,0.046875,-0.078125,0,0.015625,-0.03125,0.0078125,0.015625,-0.0078125,-0.046875,-0.0625,0.03125,-0.0390625,0.0625,0,0.015625,0.015625,0.046875,-0.0078125,-0.046875,0,0.015625,0,-0.03125,-0.0390625,0.0546875,0.046875,0.03125,0.0546875,0.0546875,0.0234375,-0.0625,-0.0390625,0.0546875,0.03125,0.046875,0.0703125,-0.0546875,0,-0.03125,0.0078125,-0.0625,-0.03125,0.0546875,0.015625,0,0.03125,0.0078125,0.0078125,-0.0390625,-0.0859375,-0.0625,0.015625,0.015625,0.0390625,0.0546875,0.03125,-0.0078125,-0.078125,0.046875,-0.09375,0.0546875,0.0078125,0.0546875,0.0625,0.0234375,-0.015625,-0.015625,0.0078125,-0.03125,-0.0703125,-0.015625,-0.046875,-0.109375,0.015625,0.015625,0,-0.0390625,0.03125,0.0625,0.0859375,-0.0234375,0.03125,-0.0234375,0.0078125,0.046875,-0.0625,-0.03125,0.046875,0.0078125,-0.015625,-0.015625,0,0,0.0078125,-0.0078125,0.0078125,0,0.03125,0.015625,0.015625,-0.046875,-0.0703125,-0.015625,-0.015625,-0.0078125,0,0.0859375,0.0078125,0.0078125,0.0625,0.0390625,-0.046875,0.0078125,0.0078125,0.015625,0.0078125,-0.046875,-0.0546875,-0.0078125,-0.0546875,-0.03125,-0.0625,-0.109375,0.125,0.1015625,-0.0078125,0,0.0078125,0.0078125,-0.0078125,-0.015625,0,-0.015625,0.0078125,-0.1015625,-0.0234375,0.0625,-0.015625,-0.046875,0.1171875,0.0546875,-0.09375,0.0546875,0.03125,-0.046875,0.046875,-0.0078125,0.09375,-0.1015625,0.0078125,0,0.0078125,0,0.0625,-0.03125,-0.0859375,0.0859375,-0.09375,-0.0859375,0.0859375,-0.0625,0.0546875,0.046875,-0.0234375,-0.0234375,-0.0078125,-0.03125,0.0234375,0.046875,0.0078125,-0.0234375,-0.0078125,-0.0390625,-0.0234375,-0.03125,-0.03125,0.015625,-0.0234375,0.046875,-0.0234375,-0.0390625,-0.03125,0.015625,0,-0.03125,0.0390625,0,0.0234375,-0.0078125,-0.015625,-0.0078125,0.0078125,0,-0.0234375,0.03125,0.015625,0.0078125,0.0078125,-0.0234375,0.015625,-0.0546875,0.015625,0.0234375,-0.046875,-0.0234375,0.03125,-0.015625,0.0078125,-0.0078125,-0.0078125,-0.1015625,-0.0546875,0.0390625,0.015625,0.0546875,-0.0234375,-0.0625,-0.03125,0.03125,-0.015625,0.0625,-0.0625,-0.046875,0.09375,-0.0078125,0,-0.015625,0,0.0078125,0,-0.0078125,0.0078125,0.0390625,0.0234375,0.0078125,-0.0546875,0.03125,0.015625,-0.0625,0.0625,-0.015625,0.0234375,0.0703125,-0.0390625,0.0234375,-0.0234375,0.0078125,-0.0546875,-0.0234375,-0.09375,0.0546875,0.0078125,0.0390625,0.0078125,0.0078125,0,-0.0234375,-0.015625,-0.0625,0.0546875,0.0859375,-0.0546875,-0.015625,-0.015625,-0.0859375,-0.078125,0.1015625,-0.0078125,0.0859375,0.0625,0.0234375,-0.078125,0.0390625,-0.078125,-0.0625,-0.0078125,0.046875,-0.015625,-0.0234375,-0.0546875,-0.03125,-0.046875,0.0078125,-0.015625,0,-0.0625,0.1015625,0.0625,-0.0703125,0.0703125,-0.015625,-0.0390625,0.0078125,0,-0.0703125,0,-0.0078125,0.015625,-0.0703125,-0.0390625,0.0546875,-0.0390625,0.015625,0.0234375,0.0390625,-0.0234375,-0.03125,0.03125,-0.0625,-0.0234375,-0.0078125,-0.015625,-0.015625,0.0859375,0.03125,-0.0546875,-0.046875,0.0234375,-0.0703125,-0.0703125,0.046875,0.0078125,0.03125,-0.0078125,-0.015625,-0.046875,-0.109375,-0.0625,0.109375,-0.015625,0.0078125,-0.046875,0.0625,-0.0234375,0.0078125,-0.046875,0,-0.0390625,0.0078125,0.0234375,-0.03125,0.0078125,-0.046875,0.0078125,-0.078125,0.0078125,0.03125,0.0625,-0.0625,0.046875,0.0390625,-0.078125,0.0625,0.015625,0.0234375,-0.0546875,-0.0078125,-0.0078125,0.03125,0.046875,-0.03125,-0.0078125,-0.0546875,0.015625,0.0546875,0.015625,-0.015625,0.0234375,-0.0234375,0.078125,0.03125,-0.0234375,-0.09375,0.0078125,-0.015625,-0.0078125,-0.015625,-0.0078125,-0.015625,-0.0078125,-0.015625,-0.0234375,0.0234375,0,-0.0078125,0,0.0078125,0.0703125,0.0078125,0.0078125,-0.0703125,-0.0390625,0.03125,-0.046875,0,0.0078125,-0.0234375,0.0078125,0.0234375,-0.046875,-0.1015625,0.046875,0.0078125,0.0234375,0.0234375,0,0.0234375,0.0234375,0.03125,0.015625,-0.0390625,0.0078125,-0.015625,0.0078125,-0.015625,0,0.015625,-0.0078125,-0.0078125,0,0,0.0078125,-0.0234375,0.0078125,0.0390625,-0.03125,-0.0234375,-0.03125,0.0078125,-0.0078125,-0.0390625,-0.046875,-0.0859375,0.0078125,0.0546875,0.0078125,-0.0390625,-0.0078125,0,0.0625,-0.03125,0.03125,0,0.046875,0,0.015625,-0.046875,-0.0546875,-0.0390625,0.0546875,-0.0234375,0,0.015625,-0.0234375,-0.03125,-0.015625,-0.015625,-0.015625,-0.0625,-0.0078125,0.0703125,-0.0390625,-0.0625,-0.0625,-0.046875,0.0078125,-0.03125,-0.015625,0.015625,0.0546875,0.0078125,-0.0546875,0.03125,-0.0078125,-0.0078125,0.0390625,-0.03125,-0.046875,-0.015625,-0.0078125,0.03125,0.015625,0,0.0390625,0.0546875,-0.0078125,0.0078125,-0.0546875,-0.015625,0.09375,-0.03125,-0.0078125,0,-0.03125,0.0546875,0.0234375,0,0.0625,-0.015625,-0.0078125,-0.03125,-0.0390625,-0.03125,0.015625,-0.0390625,-0.0234375,-0.015625,0.0625,0,-0.015625,0.0078125,0.0078125,-0.015625,0,0.0234375,0.0234375,0.0234375,0.03125,-0.0078125,0,0.0078125,-0.015625,0,0.015625,-0.0390625,0.0078125,-0.0390625,0.0390625,0.015625,-0.03125,-0.015625,0.0390625,0.1484375,0.0234375,-0.0859375,0.015625,-0.015625,0,-0.046875,-0.015625,0.03125,0.0078125,0.015625,-0.0390625,0.0390625,-0.0390625,-0.046875,-0.046875,-0.0390625,-0.0390625,0.1484375,0.015625,0.0546875,0.0625,-0.0390625,-0.0234375,0.0234375,0.1015625,0.03125,-0.0078125,-0.0390625,-0.0234375,0.0546875,-0.015625,0.0234375,0.015625,0.0390625,0.015625,0,-0.046875,0.0078125,0.0078125,0.0078125,-0.0546875,0.0078125,-0.046875,-0.0859375,0.0234375,-0.015625,0.0234375,0.046875,-0.0234375,-0.0859375,-0.0625,-0.015625,-0.015625,0.0078125,-0.046875,0.03125,0.0390625,-0.015625,-0.0703125,-0.046875,0.0234375,-0.0078125,0.0234375,0.0078125,-0.0234375,0.03125,-0.0078125,0.0234375,0.0625,-0.015625,0.0546875,0.0234375,-0.0390625,-0.0234375,-0.046875,-0.03125,0.0625,0.046875,0.0234375,-0.1171875,0.0859375,-0.046875,0.0703125,-0.015625,0.015625,0.0078125,0.0234375,-0.015625,0,0.1640625,0.03125,-0.0859375,-0.0859375,0,0.03125,-0.015625,0.0078125,0.0078125,0.0625,-0.0546875,-0.0078125,-0.109375,0.078125,0.015625,0.0078125,-0.03125,-0.015625,0,-0.0234375,-0.015625,-0.046875,-0.0078125,0.015625,0.015625,-0.03125,-0.0859375,0.015625,-0.0078125,0,0.015625,-0.0078125,0,0.0234375,-0.0234375,0.015625,-0.0078125,0.0234375,-0.0078125,0,-0.0234375,0.046875,-0.03125,0.0078125,0,-0.0078125,-0.0078125,0,0.0078125,0.015625,0,0,-0.0078125,-0.0390625,0,-0.0859375,0.0546875,-0.015625,0.0859375,-0.0234375,-0.015625,0,-0.0078125,0.0078125,-0.0234375,0.0390625,-0.0078125,0.03125,-0.0703125,-0.0625,0,-0.0078125,-0.0078125,-0.078125,-0.0078125,-0.03125,0.0859375,0.015625,0,0,0,0,0.0078125,-0.0078125,0,0,-0.015625,0,-0.015625,0,0,-0.1015625,0.015625,-0.0234375,-0.03125,-0.015625,-0.015625,0.046875,0.0078125,-0.0234375,0.1875,-0.1015625,-0.0078125,0.0546875,-0.0078125,-0.0390625,0.0390625,0.0546875,-0.015625,0.0078125,0,-0.03125,-0.0703125,-0.0234375,-0.0703125,-0.046875,0.0078125,0.0078125,0.015625,-0.0703125,-0.03125,0,-0.046875,0,0,0.0234375,-0.0078125,0,-0.0625,0,-0.0390625,-0.0625,0.0078125,-0.03125,0,0,0.078125,-0.015625,-0.0078125,-0.015625,-0.0078125,0.0078125,0.015625,-0.0078125,0,0.03125,-0.0078125,0,-0.0078125,-0.03125,-0.015625,-0.0078125,-0.0078125,0.0078125,0,-0.0390625,-0.0078125,0.015625,0,-0.015625,-0.0234375,-0.0390625,0,-0.09375,-0.140625,0,0.015625,0.03125,-0.0078125,0.0078125,0.0546875,-0.015625,-0.0078125,0.0078125,-0.046875,-0.1640625,0.046875,-0.0234375,-0.0078125,0.0078125,-0.0078125,0,0.015625,0,0.0078125,0.0078125,-0.015625,-0.015625,-0.0078125,0.015625,-0.015625,-0.03125,0.0234375,-0.015625,0.0390625,0,-0.0234375,-0.0234375,0,-0.0390625,0.03125,-0.015625,0.0859375,-0.09375,-0.046875,0,-0.0078125,0.015625,-0.015625,-0.09375,-0.0390625,0.1484375,-0.09375,0.0078125,-0.015625,-0.046875,0.0078125,-0.0234375,-0.046875,-0.0390625,0,0.03125,-0.0234375,-0.0625,-0.0234375,0.015625,-0.0546875,-0.0625,-0.015625,-0.0546875,0.03125,-0.03125,0.0078125,-0.0234375,-0.015625,-0.0625,0.0703125,-0.03125,0.015625,-0.0703125,0,0.0078125,-0.03125,0.0234375,-0.03125,-0.0390625,-0.015625,0.1015625,-0.0546875,-0.0390625,-0.046875,-0.0078125,-0.0078125,0.046875,-0.0078125,-0.015625,0.0390625,0.0390625,-0.015625,-0.0078125,0,0.0234375,-0.015625,-0.0390625,0,0,0.015625,-0.015625,-0.0078125,-0.0234375,0.0078125,0.15625,0.0078125,0,-0.03125,-0.0859375,-0.03125,-0.0078125,-0.0234375,-0.0078125,-0.046875,0.0703125,-0.0703125,0,0.03125,-0.0078125,-0.046875,-0.0703125,0,-0.0234375,0.0078125,-0.046875,-0.0234375,-0.03125,-0.0234375,-0.0078125,-0.03125,-0.0078125,0.03125,0.0625,0,-0.015625,-0.0078125,-0.015625,0.0625,-0.015625,-0.03125,0.0546875,-0.09375,-0.03125,0.0390625,-0.0078125,-0.015625,-0.0078125,-0.0078125,0.0078125,-0.078125,0.0703125,0,0.0625,-0.015625,-0.0234375,0.03125,0,0.0625,-0.0078125,-0.0078125,-0.0234375,-0.0390625,-0.1015625,-0.046875,-0.0078125,-0.015625,0.0078125,0.0078125,0.015625,0,-0.0078125,0.0234375,-0.0078125,0,-0.0078125,0.0078125,0.1015625,-0.046875,0.0546875,0.0625,-0.0859375,-0.09375,-0.0546875,-0.0234375,-0.0234375,-0.0234375,0,0.0390625,0.046875,0.03125,0.046875,-0.0078125,-0.0078125,-0.0390625,-0.0390625,0.0078125,-0.03125,-0.03125,0,0.1015625,0,0.015625,0,-0.0078125,-0.0078125,-0.0078125,-0.0078125,-0.0078125,0.0078125,-0.015625,0.0234375,-0.0703125,-0.0078125,-0.1171875,0.0703125,0.1015625,0.0390625,-0.078125,0.0859375,-0.03125,0.140625,-0.015625,-0.0625,-0.0859375,0.0703125,0.015625,0,0.0546875,0.03125,-0.0078125,0,0.015625,0.015625,-0.0078125,-0.078125,0.0234375,0.03125,-0.03125,-0.046875,0.0546875,0.0546875,-0.03125,0.0234375,-0.0703125,-0.03125,-0.015625,-0.0546875,-0.0078125,-0.0234375,-0.046875,-0.046875,-0.015625,0.109375,0.0546875,-0.0078125,-0.0546875,0,0,-0.015625,0.0390625,-0.0078125,0.0078125,0.0078125,0.0546875,0.03125,0.015625,-0.0390625,-0.0078125,-0.0078125,0,-0.0390625,-0.015625,-0.0078125,0.0078125,-0.0078125,-0.0390625,0.0078125,-0.015625,0.0859375,0.0703125,-0.03125,0.015625,-0.015625,-0.03125,-0.0546875,0.0625,-0.0703125,0.0078125,0.015625,-0.0546875,0.0078125,-0.0234375,-0.0234375,-0.0078125,0,0.03125,0.0078125,-0.0625,-0.0703125,0.015625,0.0078125,-0.0078125,-0.0078125,0.0078125,-0.015625,0,0,0.0234375,-0.03125,0.03125,0.03125,0.046875,-0.03125,-0.0078125,-0.0234375,0.0078125,-0.0078125,0.0078125,0,0.015625,-0.0390625,-0.0859375,0.046875,0.0234375,0.0234375,-0.0390625,0.0390625,0,-0.046875,0.0390625,-0.078125,0.015625,0.03125,-0.0390625,-0.0234375,0.0078125,-0.0078125,-0.03125,0.03125,0.1171875,0.0234375,-0.0625,0.0078125,-0.015625,0.0390625,-0.046875,-0.0078125,0.0234375,-0.03125,-0.015625,0,-0.015625,0.03125,0,-0.0546875,0,0.0234375,-0.0078125,0.078125,-0.046875,-0.078125,0.0078125,0.0078125,-0.046875,-0.03125,-0.140625,0,0.1015625,0.015625,-0.0859375,0.09375,-0.015625,-0.046875,-0.0234375,0.046875,-0.0078125,-0.0546875,0.0078125,-0.0390625,-0.0078125,0.03125,-0.015625,0.0390625,0,-0.0078125,-0.03125,-0.0078125,-0.0078125,-0.015625,0.09375,0.0703125,0.1015625,-0.03125,-0.03125,0,0.0546875,-0.015625,0.046875,0.015625,0.015625,-0.0390625,-0.0625,-0.0234375,-0.0546875,0.09375,0.0078125,0,-0.0390625,-0.0625,-0.0390625,-0.03125,-0.09375,-0.0078125,-0.0546875,0.078125,0.0234375,-0.0078125,0.015625,-0.0390625,0.03125,-0.0859375,0.0234375,0.078125,0.0390625,-0.0546875,-0.0078125,0.03125,-0.0390625,0.046875,-0.015625,0.0390625,-0.0703125,0.0390625,0.03125,0.0078125,0.078125,0.0703125,-0.0625,-0.0546875,-0.0390625,-0.046875,-0.1171875,0.0234375,-0.0703125,-0.015625,-0.0234375,-0.015625,0.03125,-0.0078125,0.0234375,0.0234375,0,-0.015625,-0.0078125,-0.015625,-0.015625,0.0078125,0.0078125,0,0,0.0078125,0.0390625,-0.0859375,0.0390625,0.0078125,-0.078125,0.0078125,0.0234375,-0.03125,0.0859375,0,-0.03125,0.0078125,0.0859375,-0.09375,-0.046875,0.078125,-0.078125,0.109375,-0.0703125,-0.046875,-0.0546875,-0.0625,-0.0234375,0.015625,-0.1171875,0.15625,0,0.0078125,0.0078125,-0.0078125,0.0078125,0.0078125,-0.0078125,0,0.0078125,0,-0.0390625,-0.0546875,0,-0.0078125,-0.1328125,0.1328125,0.0546875,-0.078125,0.078125,0.0625,-0.1015625,0.1171875,0.0390625,-0.1171875,-0.0078125,-0.0625,0.0625,0,-0.0234375,0.0859375,0.09375,-0.0390625,0.1640625,-0.109375,0.0390625,0.0703125,-0.0390625,0.0078125,-0.0078125,0.03125,0.0234375,-0.0234375,-0.0234375,-0.0703125,-0.0078125,-0.03125,0.0078125,0.0546875,-0.015625,0.0078125,0.0078125,0,0,-0.0234375,0.0078125,0.0078125,-0.078125,-0.0078125,-0.015625,-0.046875,0.0078125,0.015625,0.0078125,0,-0.03125,-0.0390625,-0.0078125,0.015625,-0.0625,0.0234375,0.03125,0.015625,0,-0.0234375,-0.0390625,0.0078125,-0.0703125,0.078125,-0.0625,0.03125,0.0390625,0,-0.0234375,0.046875,-0.0390625,-0.0625,-0.0390625,-0.0234375,0.0625,0,0.015625,-0.046875,0.03125,-0.046875,0.0234375,-0.03125,0.0546875,-0.09375,0.046875,-0.0390625,0.0078125,0.0078125,-0.015625,-0.015625,0,-0.03125,-0.015625,0.015625,0.0234375,0.0390625,-0.0234375,0.046875,0.0234375,0.03125,-0.0078125,0.0546875,0,0.0625,0.09375,-0.0390625,0.0625,-0.0078125,-0.0234375,-0.0859375,0.0078125,-0.0390625,-0.0234375,0.0234375,-0.015625,0.0234375,-0.03125,0.03125,-0.0625,-0.015625,0.03125,-0.0390625,0,-0.0703125,0.015625,-0.015625,-0.0390625,-0.0546875,-0.0546875,0.0234375,0.0234375,-0.015625,-0.0859375,0.0078125,-0.0703125,-0.0703125,0.046875,-0.15625,0.1875,-0.09375,0.0234375,-0.0234375,-0.0078125,0.0625,0.046875,-0.0390625,0.0859375,-0.078125,0.03125,0.0625,0.015625,0.03125,0,-0.0078125,-0.078125,-0.0390625,-0.0625,0.0234375,-0.0703125,0.046875,0.0390625,-0.0703125,0.0546875,0.0390625,0.078125,0.0078125,0.109375,0.015625,0.078125,0.0234375,0.015625,-0.0703125,-0.015625,-0.03125,0.078125,-0.0078125,0.0234375,-0.0234375,0,0,0.046875,0.015625,-0.0703125,0.140625,0,0.015625,0.0703125,0.046875,-0.015625,0.0390625,-0.0234375,-0.0234375,-0.0625,-0.0234375,-0.0390625,-0.03125,-0.0859375,-0.0703125,-0.046875,-0.0234375,-0.09375,0.03125,0,0.015625,-0.0546875,-0.0078125,-0.046875,-0.140625,-0.1171875,-0.0078125,0.015625,-0.0234375,-0.03125,-0.140625,-0.015625,0.015625,-0.0390625,-0.0546875,-0.015625,-0.046875,0.0703125,0.0859375,0.0234375,0.0078125,-0.0625,-0.0390625,0.0390625,0.03125,0.0546875,-0.0234375,0.0078125,0.203125,0,-0.1015625,0.03125,-0.0390625,-0.0546875,-0.0546875,0,0.015625,-0.0078125,0.0078125,0.0078125,0.015625,-0.0234375,-0.0078125,0.0078125,0,0.0546875,0.0390625,-0.0078125,-0.078125,-0.1015625,-0.0546875,0,-0.0703125,0.03125,-0.046875,-0.015625,0.0703125,0.0625,-0.046875,0.0078125,0.0078125,-0.0390625,0,-0.046875,-0.0625,-0.0625,-0.03125,0.046875,-0.046875,-0.0078125,0.0078125,-0.0078125,0.015625,-0.0078125,0.0078125,-0.0078125,0.0078125,0.0078125,0.0078125,-0.0078125,0,-0.0703125,-0.0390625,0.0234375,-0.0546875,0.0234375,-0.0234375,-0.0703125,0,-0.0703125,-0.03125,-0.0390625,-0.046875,-0.09375,0.015625,0.046875,0.0546875,0.046875,0.0078125,0.09375,-0.0078125,0.03125,0.03125,-0.0859375,0.015625,-0.046875,-0.0625,0.0078125,-0.0078125,-0.078125,-0.0078125,-0.046875,0.03125,0.0078125,-0.0390625,0.0234375,0.015625,-0.015625,0.0859375,-0.0078125,-0.0078125,0.0078125,0.1171875,0.015625,-0.0390625,0.0078125,0,-0.015625,-0.0078125,-0.0234375,-0.015625,-0.0625,-0.046875,-0.015625,-0.0546875,0.0234375,-0.0234375,0.0234375,-0.0234375,-0.0546875,0.0078125,0.015625,0.0078125,0.0078125,-0.0234375,-0.03125,0.015625,0.0078125,-0.046875,-0.0390625,0.0078125,0.03125,-0.0546875,0.015625,-0.046875,0.03125,-0.1171875,0.046875,-0.0625,-0.015625,0.015625,0.03125,0.0703125,0.0078125,-0.046875,0.09375,-0.046875,0.03125,-0.03125,-0.015625,0.0859375,-0.0078125,-0.0234375,0,0.03125,0.0390625,0,0.03125,0.015625,0.0078125,-0.015625,-0.015625,-0.0234375,-0.0625,-0.0078125,-0.03125,-0.015625,-0.0078125,0.0234375,0.0546875,0.0546875,0.03125,0.0234375,-0.03125,-0.078125,0.0390625,0.078125,0.03125,-0.0078125,0.015625,0,-0.109375,0.046875,-0.078125,-0.0859375,-0.0546875,-0.046875,0.0546875,0.0234375,0.0703125,-0.09375,0.109375,-0.1171875,0.03125,-0.0390625,-0.0078125,0.015625,-0.0546875,0.0234375,0.0390625,-0.0078125,0.0703125,0.0546875,-0.078125,0.0546875,0.03125,0.0078125,0.0703125,0,-0.03125,0.015625,-0.0078125,-0.046875,0.015625,0.09375,-0.0390625,0.0390625,-0.0390625,-0.1171875,-0.0859375,0.0078125,0.0859375,0.0546875,0.0390625,0.0390625,-0.0078125,-0.0078125,0.0703125,-0.0625,0,-0.046875,0.0234375,0.0625,-0.0234375,0.046875,0.015625,0.015625,-0.0546875,0.0234375,0.046875,0.0078125,-0.0078125,-0.0234375,-0.0078125,0.0078125,-0.015625,-0.015625,-0.0234375,0.0078125,-0.03125,0.015625,-0.046875,0.0625,-0.03125,-0.015625,0.046875,-0.0546875,-0.1328125,-0.0078125,0,-0.1171875,-0.0546875,-0.015625,0,-0.0546875,0.0625,0.1796875,0.0078125,0,0,0.03125,0,-0.0546875,0.09375,-0.0703125,0.0390625,-0.0390625,0.03125,0.015625,0.046875,-0.0703125,0,-0.046875,0.046875,0.0390625,0.0703125,0.078125,-0.03125,0.046875,0,-0.0703125,0.0390625,-0.1015625,-0.0625,-0.0234375,0.0546875,-0.0234375,-0.0390625,0.0234375,0.015625,0.0234375,-0.015625,0,-0.015625,-0.015625,0.0078125,-0.015625,0,0,-0.0078125,-0.015625,0,0,-0.0234375,-0.015625,0.015625,-0.0546875,-0.0390625,-0.0703125,0.109375,-0.03125,-0.0546875,-0.03125,-0.0546875,-0.03125,0.0234375,-0.0390625,-0.015625,0.015625,0.03125,-0.015625,0.015625,-0.03125,-0.03125,0.0546875,0,0.0625,0.046875,-0.0625,-0.015625,0,0,0.0078125,0,-0.0078125,0.015625,-0.0078125,0,-0.0078125,-0.0546875,-0.046875,-0.0546875,-0.015625,-0.1015625,0.0625,0.0625,-0.0859375,0.078125,-0.0546875,-0.015625,0.0078125,0,0.0390625,-0.0078125,-0.0703125,0.015625,0.015625,0.0234375,-0.046875,-0.0078125,0.1328125,0.0625,0.0703125,0.015625,-0.125,-0.0625,0.0234375,0,0.015625,0.015625,0.0390625,-0.0234375,0.0703125,0.0546875,-0.03125,0.0078125,0.0234375,0.015625,0.03125,-0.0234375,-0.0390625,-0.0234375,-0.0390625,0.0546875,0.015625,-0.0234375,-0.0234375,-0.0234375,-0.0625,-0.046875,-0.0234375,-0.0390625,0.0078125,-0.0078125,-0.015625,-0.03125,0.015625,0,-0.0078125,0.0078125,0.015625,0,0,-0.0234375,0,-0.015625,0.0078125,0.0078125,-0.046875,-0.0625,-0.03125,0.0390625,0.1015625,-0.0546875,0,-0.0546875,-0.0703125,-0.0546875,0.0390625,0.0234375,0.0078125,0,-0.046875,-0.0234375,0,0.0625,-0.0078125,-0.0078125,0.0390625,0,0,-0.0234375,0,-0.015625,0,-0.015625,-0.015625,-0.0078125,0.0546875,0,0.0234375,0.0078125,0.046875,-0.0546875,0.0078125,0.0078125,-0.0078125,-0.0234375,0.0546875,-0.1015625,0.03125,-0.015625,-0.03125,-0.015625,0.0390625,-0.03125,-0.0625,-0.015625,-0.015625,-0.0234375,0.0390625,-0.0078125,-0.03125,0.109375,0.0546875,-0.0234375,0.0390625,-0.03125,-0.0390625,-0.1015625,0.0078125,0.0078125,-0.015625,0.0078125,-0.0546875,-0.015625,-0.03125,0.015625,0.0390625,-0.03125,0.0703125,-0.0234375,0.0546875,-0.015625,0.109375,-0.046875,-0.0703125,-0.0625,0,0.0078125,0,-0.0546875,0.0390625,-0.015625,-0.0625,-0.1015625,0.078125,-0.0234375,-0.0546875,0.015625,-0.046875,0.0859375,0.0078125,0.046875,0.015625,0.03125,0.0234375,0.0234375,-0.0546875,-0.0078125,-0.015625,0.015625,0.0390625,-0.0546875,-0.046875,0.0078125,-0.015625,0.0390625,0.0390625,0.015625,-0.046875,-0.0234375,0.0078125,-0.0234375,-0.015625,0.015625,-0.0078125,-0.0078125,0,-0.03125,0.0390625,-0.015625,0,-0.0546875,-0.0546875,-0.046875,0.0078125,-0.09375,0.0390625,-0.0078125,0.015625,0.0234375,0.0546875,0.046875,-0.03125,0.0234375,-0.0703125,0.1171875,0.0078125,-0.046875,-0.078125,-0.015625,-0.03125,-0.015625,0.0390625,-0.015625,0.0234375,-0.03125,-0.03125,-0.0234375,0.0390625,0.015625,0.015625,-0.0234375,-0.03125,0.03125,-0.0625,-0.0546875,0.0234375,-0.0546875,0.03125,-0.0546875,0.0078125,0.0390625,0.125,-0.015625,0.0078125,-0.0078125,0.03125,-0.0859375,-0.0390625,-0.0078125,0.015625,-0.0078125,0,-0.015625,0.0078125,0.0078125,-0.0078125,0.015625,0,0.078125,0.0859375,0,-0.0859375,-0.0703125,-0.0390625,-0.0234375,-0.03125,0.0078125,0.0234375,0.0234375,0.0703125,-0.0625,0.015625,-0.0859375,0.0625,0.015625,0.0546875,-0.0078125,-0.0234375,0.046875,0,-0.0390625,-0.015625,-0.015625,-0.0234375,0.0078125,-0.0078125,0.0234375,0.0078125,0,-0.0078125,0,0,0.015625,0.0078125,0.0703125,-0.0625,0.078125,0,-0.0234375,0.109375,0.03125,-0.0078125,0.0390625,-0.03125,-0.0546875,-0.03125,-0.0390625,0.03125,-0.0625,0.0078125,0.0078125,0.0390625,-0.0078125,-0.015625,-0.0078125,-0.015625,0.0546875,-0.0625,0.0625,0.109375,0.0390625,0.0234375,0.0390625,0,-0.0546875,-0.0546875,0.0625,0.0234375,0.0078125,0.0234375,-0.03125,-0.015625,-0.0546875,-0.015625,0,-0.046875,-0.0234375,-0.1484375,-0.0078125,0.0078125,-0.0234375,-0.0546875,0,0.015625,-0.0078125,-0.0078125,0.015625,-0.0390625,-0.015625,-0.0546875,-0.0390625,0.015625,0.0546875,0.0078125,0,0.0078125,0.0390625,-0.0234375,0.0078125,-0.03125,-0.0625,0.0078125,-0.0390625,-0.03125,0.015625,-0.0078125,-0.046875,0.0234375,-0.0625,0.0625,-0.078125,-0.0234375,0.0078125,-0.0390625,0.015625,-0.0546875,-0.0234375,-0.03125,0.046875,0,0.0703125,-0.0078125,0.03125,-0.03125,0,0,0.0078125,0,-0.0078125,0,0.0234375,0.03125,0.0234375,0.015625,-0.015625,-0.0703125,-0.0625,-0.0625,0.015625,0.0390625,-0.0078125,0.0078125,0.046875,0,0.046875,0.03125,-0.015625,0.046875,-0.0234375,-0.0390625,0.015625,0,0.015625,0,0.03125,-0.0546875,0.015625,0.0546875,-0.0546875,0.015625,-0.0625,0.046875,-0.015625,-0.09375,0.0078125,-0.1015625,0.03125,-0.015625,0.046875,0,-0.0390625,-0.1171875,0.0390625,-0.078125,0.0234375,0.0234375,0,0.015625,0.03125,0.0859375,0.0546875,-0.0859375,-0.0625,-0.0234375,0.0078125,-0.0625,0.0546875,0.015625,-0.046875,0.0390625,-0.03125,0.03125,-0.0234375,-0.0078125,0.046875,-0.0078125,0,0.0078125,-0.0078125,-0.0234375,-0.03125,0.015625,-0.0234375,0.046875,0.0390625,-0.078125,-0.0078125,-0.03125,-0.0078125,0.015625,-0.0859375,0.0234375,0.0859375,0,0.03125,-0.0390625,0,0.03125,-0.0390625,-0.015625,0.03125,0.09375,0.03125,-0.0703125,-0.0625,-0.0078125,0.0546875,0.0546875,0.015625,0,0.109375,-0.0390625,-0.078125,0.0703125,-0.046875,0.0625,0.0234375,-0.0703125,-0.03125,-0.0859375,0.0078125,0,0,0.03125,-0.015625,-0.140625,-0.0625,0.09375,-0.140625,0.1328125,-0.0234375,0.0234375,-0.0078125,-0.0703125,-0.0078125,0.0234375,-0.0234375,0.015625,0.078125,-0.0078125,0.03125,0.0078125,0.0703125,-0.078125,0.0390625,0.0078125,0,-0.078125,0.0390625,0.125,0.0546875,-0.0234375,-0.0390625,0,0.046875,-0.03125,-0.0390625,0.0078125,0.0078125,-0.0078125,-0.0078125,0.0078125,-0.015625,-0.0078125,-0.0078125,-0.015625,-0.0703125,-0.015625,0.03125,0.0703125,-0.0390625,-0.015625,-0.015625,0.0078125,-0.0234375,-0.015625,0.0078125,-0.0234375,-0.015625,0.015625,-0.0078125,0.0078125,0.0078125,-0.03125,-0.0078125,0.015625,-0.0234375,-0.0390625,-0.0625,-0.03125,0.0234375,0.015625,-0.0390625,-0.0078125,0.0234375,0,-0.0078125,0.0078125,0.015625,-0.0078125,-0.0078125,-0.0078125,0.03125,0.046875,-0.03125,-0.0234375,0.0390625,-0.0625,0.046875,0,-0.0390625,0,0.078125,-0.0546875,-0.015625,-0.0546875,-0.0703125,0.015625,0.0234375,-0.0234375,0.015625,0.0234375,-0.0078125,-0.046875,-0.0078125,-0.03125,0.0390625,0.0703125,-0.015625,-0.0078125,0,0.0546875,0.0234375,-0.015625,0.03125,0,0,-0.0078125,0.0078125,-0.0234375,0.0234375,0.0078125,-0.0625,-0.0390625,0.0703125,-0.0078125,-0.03125,-0.015625,0.0078125,-0.0078125,-0.0234375,-0.0234375,-0.0234375,-0.015625,-0.015625,-0.03125,-0.0078125,0.0078125,-0.015625,-0.015625,-0.015625,-0.0078125,0.0234375,0,-0.0078125,-0.0078125,0,-0.0078125,-0.0234375,0.015625,0,0.0234375,0,0.03125,-0.0625,-0.0703125,0.0546875,0.0859375,-0.0234375,0.0859375,0.078125,0.0234375,-0.0078125,0.03125,0.015625,-0.0625,-0.0625,0.0390625,-0.0078125,0.046875,0.0390625,-0.0390625,0,0,0,0,0.0078125,0,-0.03125,0.0234375,0.0234375,0.015625,0.015625,0.0078125,-0.015625,-0.0078125,-0.0234375,0,-0.0234375,-0.0078125,-0.0234375,-0.0546875,-0.0390625,0,-0.015625,0.03125,0.015625,0,0,0.0078125,0.0234375,0.109375,0.0546875,-0.046875,0,0.03125,-0.0546875,-0.03125,-0.0625,-0.0625,-0.015625,-0.0234375,-0.015625,-0.0625,-0.0546875,0.1015625,0.0546875,0.0390625,-0.0078125,0.015625,-0.03125,-0.0390625,-0.0625,-0.046875,0.0546875,0.0234375,-0.03125,-0.0078125,0.0078125,-0.0546875,0,-0.0234375,-0.0078125,0.0234375,-0.0390625,-0.0390625,-0.03125,0.0703125,-0.0546875,0.0625,0.0703125,-0.0625,-0.03125,-0.078125,0.015625,0.015625,0.015625,0.0390625,-0.0078125,-0.015625,-0.0390625,-0.03125,-0.0234375,0,-0.046875,-0.03125,-0.015625,-0.0546875,-0.046875,0.03125,0.015625,0.015625,-0.0625,0.015625,-0.0546875,-0.0234375,-0.0078125,-0.0703125,0.0078125,0.0078125,-0.0078125,-0.0078125,-0.0078125,-0.03125,0.125,-0.0625,0.0390625,-0.0078125,-0.046875,0.0390625,-0.046875,0.0625,0.1015625,-0.03125,-0.03125,-0.015625,-0.0625,0.046875,0,0.0234375,-0.0546875,0.0234375,-0.046875,0,0.0078125,0.0078125,-0.0234375,0.015625,-0.0078125,-0.0234375,-0.03125,-0.015625,-0.03125,-0.015625,0.0078125,0.0390625,-0.0234375,0.09375,0.078125,0.078125,-0.046875,-0.0390625,-0.03125,0.03125,0.0078125,-0.015625,0.0703125,0.0546875,0.015625,-0.0078125,0.203125,-0.0546875,0.0078125,-0.0078125,-0.03125,-0.0078125,-0.0078125,0.015625,0.0078125,0,0,-0.0078125,0.0078125,-0.0078125,0.03125,-0.0546875,-0.0390625,0.0703125,-0.0078125,-0.03125,-0.0234375,-0.0234375,-0.0625,-0.0078125,0.0390625,0.0078125,0.046875,0.046875,-0.0078125,0.0625,0.0078125,-0.015625,-0.0390625,-0.0234375,-0.0703125,-0.0390625,-0.0078125,-0.03125,0.015625,0,-0.0625,0.015625,-0.0078125,-0.0078125,0,0.015625,-0.0078125,0,0.0078125,0,-0.0390625,-0.015625,-0.046875,-0.0078125,-0.03125,-0.015625,0.0390625,-0.0078125,0.015625,0.0703125,-0.0390625,0.09375,-0.046875,0.0234375,-0.078125,-0.0078125,-0.0078125,-0.0234375,0.046875,0.03125,0.0234375,0,-0.046875,-0.03125,-0.0234375,-0.1171875,0.0078125,0.0625,-0.0546875,-0.015625,-0.03125,0.0234375,-0.015625,-0.0703125,-0.0234375,0,-0.078125,0.0234375,-0.0703125,-0.0234375,0.0234375,0,0.1328125,-0.015625,0.1484375,0,0.0078125,0.03125,-0.03125,-0.046875,-0.046875,-0.015625,-0.015625,-0.0390625,0.046875,-0.0234375,0.015625,-0.015625,-0.0625,0.0078125,-0.015625,-0.0078125,0.0390625,-0.0078125,-0.0078125,0.0234375,-0.046875,-0.0390625,-0.03125,0.0390625,0.015625,-0.015625,-0.015625,0,-0.015625,-0.046875,0.0703125,-0.0546875,0.03125,-0.046875,0.015625,0,-0.078125,-0.078125,0.0078125,-0.046875,0.0390625,0.015625,-0.0078125,0.0390625,0.015625,0,0.0078125,0,-0.0078125,-0.0234375,0.015625,0.0234375,-0.0078125,0.0390625,0,-0.015625,-0.0390625,-0.0234375,-0.0546875,0.015625,0.0078125,-0.0390625,0.015625,0.046875,0.0234375,0.046875,0.0390625,-0.0703125,-0.0078125,0.046875,-0.0390625,-0.0078125,0.03125,0.015625,-0.0546875,0.0234375,-0.046875,-0.109375,-0.0390625,-0.0546875,0.0078125,-0.0859375,-0.015625,0.0078125,-0.015625,-0.0234375,-0.0859375,0.0078125,-0.046875,0.015625,-0.0078125,0,-0.0078125,-0.03125,0.03125,0.0546875,-0.0703125,0.0625,0.015625,0,0.0703125,0.0234375,-0.0703125,-0.0390625,0,0,-0.03125,0.078125,-0.0625,0,0.046875,-0.125,0.0546875,0.0078125,0,-0.0625,0.015625,0.0078125,0,-0.046875,-0.03125,0,0.015625,-0.078125,-0.03125,0.0625,-0.03125,0.1171875,0,-0.0390625,0.0546875,-0.0546875,-0.0390625,-0.03125,0.03125,0.0078125,0.015625,0.0078125,-0.015625,-0.0546875,-0.0703125,-0.03125,-0.046875,0.046875,-0.1171875,0,0.0859375,-0.0390625,0.0859375,-0.046875,-0.1015625,0.03125,-0.0546875,-0.0546875,-0.0078125,-0.015625,-0.0625,-0.0546875,0.0390625,0.1171875,0.078125,0.0546875,-0.03125,0.0234375,-0.0625,-0.0390625,0.015625,-0.03125,0.0859375,0.109375,-0.0078125,-0.0234375,0.0625,-0.046875,0.03125,0.015625,-0.0625,0,-0.0234375,0.0546875,-0.0625,0.015625,0.0546875,0.03125,0.0625,0.0234375,-0.046875,0.015625,-0.0078125,-0.0859375,-0.015625,-0.0078125,0.015625,0.0859375,0.03125,-0.0078125,0.0234375,0.015625,-0.0078125,-0.0078125,0,0.015625,-0.015625,-0.0078125,-0.0078125,-0.015625,-0.03125,-0.0234375,-0.0390625,0.0625,-0.078125,0.046875,0.0390625,-0.0078125,0.046875,-0.0078125,-0.0078125,0.0546875,-0.0078125,-0.0625,-0.0234375,0.0703125,-0.0390625,0.0390625,-0.0390625,0.0078125,0,-0.03125,0.0859375,0.0546875,-0.015625,-0.015625,-0.0625,0,-0.0078125,0,0.0078125,-0.0078125,-0.0078125,0.0078125,0.0078125,0.0078125,-0.015625,-0.0234375,-0.0078125,0.0546875,0.03125,-0.015625,0,0.0390625,-0.0625,-0.015625,-0.0234375,-0.0234375,0.1015625,-0.015625,0.15625,0.0546875,-0.0625,0.0234375,0.0234375,0,0.0078125,-0.0703125,-0.03125,0,-0.046875,-0.0234375,0.046875,0.0078125,0.03125,0.0078125,0.015625,0,0.0078125,-0.0078125,-0.0078125,0.015625,-0.0234375,-0.0859375,-0.0234375,0,-0.09375,0.046875,0.015625,0.015625,0,-0.0234375,-0.0390625,-0.0078125,0,-0.0390625,-0.0234375,0,-0.015625,0.015625,0,-0.03125,-0.03125,0.0625,-0.0078125,0.0546875,0.0078125,0,0.0390625,0.015625,0.0078125,-0.0078125,0.03125,0.03125,-0.046875,-0.03125,0,-0.0234375,-0.03125,-0.0234375,0.0078125,-0.0390625,0.03125,-0.0390625,0.046875,-0.046875,0.0078125,0.0078125,0.015625,-0.0078125,-0.0234375,0.1015625,0.0859375,0,0.0390625,-0.0234375,0,-0.0078125,0,-0.0078125,-0.015625,-0.015625,0.0078125,0,0,-0.015625,0.0078125,-0.046875,0.0234375,-0.0546875,-0.0625,0.0078125,-0.03125,-0.0078125,-0.03125,0.0234375,0.03125,-0.03125,0.0078125,-0.015625,-0.0078125,-0.03125,0,0,0,0.046875,-0.03125,0.0546875,-0.0234375,-0.0390625,-0.1328125,-0.0390625,-0.015625,-0.0546875,0.0234375,0.0234375,0.078125,0.046875,0.015625,-0.0078125,-0.0078125,-0.0078125,-0.03125,0.1015625,0.046875,0.0390625,0.0078125,-0.0390625,-0.078125,-0.0625,-0.0234375,-0.03125,-0.0390625,0.0546875,-0.0078125,0.0078125,-0.0234375,-0.03125,0.0703125,-0.0390625,-0.015625,-0.0078125,-0.09375,0.0234375,-0.0546875,0.046875,0.0078125,-0.0390625,-0.0234375,-0.0078125,-0.015625,-0.046875,-0.046875,-0.046875,-0.015625,-0.0234375,0.015625,-0.0078125,0.015625,0.0234375,-0.0546875,-0.1328125,-0.0625,-0.078125,-0.0546875,-0.0625,-0.0234375,-0.03125,0.015625,0.0546875,0.0390625,0.015625,0.0078125,0.046875,0.0546875,-0.046875,0.0546875,-0.015625,0.0390625,-0.015625,-0.078125,-0.03125,-0.0703125,-0.1171875,0.015625,-0.0234375,0.0078125,-0.0703125,0.0546875,0,-0.0234375,0.0234375,-0.0625,-0.03125,0.09375,-0.0078125,-0.0234375,-0.1015625,0,0.0234375,-0.03125,-0.015625,0.015625,-0.0234375,-0.0390625,0.03125,0.0390625,0.0859375,-0.015625,0.03125,-0.0078125,-0.0234375,0.03125,-0.015625,-0.078125,-0.046875,-0.03125,0,-0.03125,-0.0234375,0.0390625,0.0078125,0.03125,0,-0.0078125,0.09375,0.0078125,0,-0.046875,-0.015625,0.0078125,0,0.0078125,-0.0078125,-0.015625,0,0,-0.0078125,-0.015625,0.03125,0.0078125,-0.0234375,0,0.015625,0.0078125,0.0234375,-0.0078125,0.046875,-0.0546875,-0.03125,0.0546875,0.0078125,-0.0234375,0.015625,-0.015625,0,0.03125,0.1640625,-0.0390625,0.0546875,0.0078125,-0.078125,-0.0703125,-0.0234375,-0.015625,0,-0.0078125,0.015625,0.0078125,-0.0078125,0.015625,0,0.0078125,0.015625,0.0390625,0.0625,0.015625,-0.015625,-0.0625,-0.1015625,-0.03125,0.03125,0.015625,0.0234375,0.078125,-0.0078125,-0.015625,0.015625,0.0390625,0.0390625,-0.0078125,-0.03125,-0.0703125,0.125,0.015625,0,-0.03125,-0.0390625,0.0078125,-0.03125,0.0390625,0.0234375,0.0078125,-0.015625,0.015625,0.03125,0.03125,-0.0234375,0.0078125,-0.0078125,-0.0390625,0.015625,0,0.0703125,0.0703125,-0.03125,-0.0234375,-0.03125,-0.0078125,0.0390625,0.0078125,-0.046875,-0.03125,-0.03125,-0.0546875,-0.0390625,-0.03125,-0.0234375,-0.0078125,0.0078125,0.0078125,-0.0078125,0,0,0,0.0078125,-0.015625,-0.0234375,0.0234375,0.0234375,-0.046875,-0.078125,-0.015625,0.015625,0.015625,0.0546875,-0.03125,0.015625,0.0546875,0.0703125,-0.1015625,-0.03125,0.046875,-0.0078125,0.015625,-0.0390625,0.03125,0.046875,-0.1015625,-0.078125,0.015625,0.0234375,0.03125,0,0.0078125,-0.0078125,0,0,0.0078125,0,0,0,-0.015625,0.0234375,-0.046875,0.0234375,0.0078125,0,-0.0234375,-0.03125,-0.0390625,-0.03125,-0.0625,-0.0546875,-0.03125,-0.0234375,0.03125,0.0234375,-0.0546875,0.015625,-0.046875,-0.0390625,0.09375,-0.0234375,0.0078125,0.0703125,-0.0859375,0.0390625,0.0234375,-0.015625,0,-0.03125,-0.0234375,-0.0859375,-0.03125,-0.078125,-0.0078125,0.0234375,0.0078125,0.078125,0,0.0390625,-0.0078125,-0.0390625,0.015625,-0.0078125,-0.0234375,0.0234375,0.0234375,0.09375,0.0234375,-0.03125,0.0390625,-0.015625,-0.015625,0.03125,-0.015625,-0.0078125,-0.0546875,-0.046875,0.0234375,0,0,-0.0390625,-0.0078125,-0.03125,0.0703125,-0.0390625,0.03125,0.015625,0,-0.078125,-0.0625,-0.0234375,0,0.015625,0.0703125,0,-0.03125,-0.0625,0,-0.078125,0,-0.046875,-0.046875,0.0546875,0.0546875,-0.0546875,0.0625,0,-0.0078125,-0.0390625,0.0078125,0.0078125,0.0078125,0.0078125,-0.0703125,-0.125,-0.0234375,-0.0234375,-0.0234375,0.0703125,-0.0078125,0,-0.0703125,0.125,-0.0234375,0.0078125,-0.0234375,0.0234375,0,-0.0546875,0.0078125,-0.046875,-0.0078125,-0.0390625,0.046875,-0.0546875,0.03125,-0.0078125,-0.0625,0.125,0.03125,-0.0234375,0.03125,0.015625,0.0078125,0.015625,-0.0234375,0.0078125,-0.0234375,0.0078125,-0.046875,0.015625,0.0546875,-0.015625,-0.0546875,-0.0546875,-0.03125,-0.03125,-0.03125,-0.03125,0.0546875,-0.0078125,-0.0390625,-0.0234375,-0.015625,0,-0.015625,-0.0078125,-0.0078125,0.0078125,0,0.015625,0.015625,0,-0.015625,0.0078125,-0.0234375,0.0078125,-0.0390625,-0.0390625,-0.046875,-0.0390625,0.0078125,0.03125,-0.03125,0.0390625,0,0.0078125,-0.0078125,-0.03125,0.0078125,-0.015625,0.0625,0.078125,-0.0625,-0.0703125,-0.0390625,-0.0234375,0,-0.03125,0,0.0078125,0,-0.0078125,-0.0078125,0,0.0078125,0,0,0.0078125,0.0234375,0.0078125,0.0546875,-0.0234375,0,-0.0234375,0.0546875,-0.03125,-0.0390625,0.03125,-0.0078125,-0.0078125,-0.0703125,-0.0078125,-0.0390625,0.0078125,0.0234375,0,-0.0390625,-0.0078125,0.0078125,0.0390625,0.09375,-0.0546875,0,-0.015625,-0.03125,-0.0078125,-0.0390625,-0.03125,0.078125,0.015625,0.0078125,-0.015625,0.0078125,0.0390625,-0.0546875,-0.0234375,0.03125,-0.0703125,-0.0234375,0.0078125,-0.0234375,0,-0.015625,0,0.015625,0.0078125,-0.015625,0.0078125,0,0.015625,0.0234375,-0.015625,-0.0078125,0,0.015625,0.015625,0.0078125,-0.0234375,0,0.0078125,0.0078125,0.0078125,-0.0078125,0,0.0390625,0,-0.03125,0,-0.046875,0,-0.0390625,0.015625,-0.0078125,-0.0078125,0.109375,0,-0.046875,-0.0234375,-0.0390625,-0.015625,-0.015625,-0.015625,0.0078125,0.03125,-0.03125,0.015625,-0.0078125,-0.0078125,0,0.015625,0,-0.015625,-0.015625,-0.015625,0.0078125,0.0078125,0.0078125,0.015625,-0.0234375,0.03125,0,0,-0.03125,-0.0234375,0.0078125,-0.0078125,0.0546875,0.0078125,0,0.015625,-0.0546875,-0.015625,-0.0078125,0,0.0078125,0.0078125,0.03125,-0.0078125,0.0234375,0.0546875,0.03125,-0.0390625,-0.015625,-0.0234375,0.0703125,0,-0.03125,-0.0625,-0.0703125,-0.046875,0.0625,0,-0.0234375,-0.0234375,-0.0234375,0,0.0234375,-0.046875,-0.03125,-0.0390625,-0.0234375,0.0234375,-0.015625,-0.0078125,-0.03125,-0.0234375,0.0078125,-0.0078125,-0.015625,0.0078125,0,0.046875,0.015625,0,0.078125,-0.03125,-0.046875,0.0078125,-0.015625,0.0234375,-0.0390625,0,-0.0078125,0.015625,0.0078125,-0.0078125,-0.03125,-0.0078125,-0.015625,-0.0078125,0.046875,0.015625,0.0625,0.0078125,0,0.0234375,-0.015625,0,-0.046875,-0.046875,0,-0.09375,-0.0859375,-0.03125,-0.0390625,0.0078125,0,0.09375,-0.046875,-0.046875,0.1171875,-0.0546875,0.0234375,-0.0234375,-0.046875,-0.015625,0.0078125,0.078125,0.015625,-0.09375,-0.0078125,-0.015625,0,0.0078125,0.015625,-0.015625,-0.03125,-0.0078125,-0.0234375,0.015625,0.0234375,-0.03125,-0.0703125,0.0625,-0.03125,0.0859375,-0.0078125,-0.0078125,0.0234375,0,0.0390625,0.0078125,0.015625,0.015625,-0.0078125,0,0.078125,-0.1015625,0.015625,0,0,0.0390625,0.0546875,-0.0625,0.0078125,-0.0625,-0.015625,0,-0.0234375,-0.0625,0.125,0.0078125,-0.0078125,-0.0078125,0.0234375,0,0,-0.0078125,0.0078125,0.015625,-0.0234375,-0.0234375,0.0078125,0.0078125,-0.046875,0.140625,0.0234375,-0.046875,-0.015625,-0.0078125,0.0390625,0,-0.015625,-0.0546875,0.078125,0.0234375,0.015625,-0.0078125,0.03125,0.0859375,-0.015625,-0.0234375,-0.0625,-0.03125,-0.0390625,0.03125,-0.015625,0.015625,-0.0078125,0.0078125,0.0078125,0.0078125,0.015625,-0.015625,-0.0078125,0,0.0234375,0.0078125,-0.0390625,0,0.0390625,-0.03125,0.03125,-0.0625,0.0078125,-0.0234375,-0.0234375,0.03125,0,-0.0234375,0.0078125,0.015625,-0.0390625,0.015625,0.0546875,0,-0.0546875,-0.0859375,-0.046875,-0.046875,0,-0.046875,0.03125,-0.046875,-0.046875,-0.0390625,0.0078125,-0.015625,-0.0390625,0.03125,-0.03125,-0.0078125,0.046875,-0.046875,-0.0078125,0.0078125,-0.03125,-0.015625,-0.0859375,0.03125,0.046875,-0.0078125,0.0625,0.0078125,0.0390625,0.015625,-0.015625,0.0078125,0.0078125,0.015625,0,-0.015625,-0.015625,0.0078125,0.03125,0.0078125,-0.015625,0.015625,-0.015625,0.0234375,0.0078125,0.015625,-0.0234375,-0.0078125,-0.0234375,-0.03125,-0.015625,-0.0234375,0.1171875,-0.0625,-0.03125,-0.0234375,-0.0234375,-0.03125,-0.046875,-0.015625,0.0546875,0.0390625,0.0078125,-0.0234375,-0.0234375,0,0.03125,-0.0390625,0,0,-0.015625,-0.0078125,0.0078125,-0.0078125,0.0234375,0.0234375,-0.0078125,0,-0.0078125,-0.015625,-0.03125,-0.015625,0.03125,-0.0078125,0,0.0234375,0,0.015625,-0.0078125,-0.0234375,0,-0.03125,0.0078125,-0.0078125,-0.046875,0.015625,-0.0078125,-0.0078125,-0.0390625,0,0.0078125,-0.015625,0,-0.03125,0.0390625,-0.015625,0.03125,-0.0546875,0.015625,-0.0234375,0,0.0078125,-0.0390625,0.046875,0.0625,0.0234375,0.0078125,-0.0234375,0.0390625,0.03125,-0.046875,-0.0625,-0.0234375,-0.046875,-0.0625,-0.046875,0,0.0703125,0.015625,0.046875,0.046875,-0.0234375,-0.015625,0.0625,0,0.078125,-0.015625,-0.1171875,-0.0859375,-0.0078125,0.0234375,-0.0390625,-0.0390625,0,-0.0234375,0.0625,-0.046875,0,-0.0390625,0.015625,0.0234375,0.03125,0.0078125,-0.015625,0.0703125,0,-0.0078125,0.0546875,0.0390625,-0.0390625,-0.0234375,0.0546875,0.0703125,-0.0703125,0.078125,0.0546875,-0.015625,-0.015625,-0.0546875,-0.03125,-0.0078125,0.0078125,-0.046875,-0.0625,-0.0078125,0.015625,0.03125,-0.03125,0.0078125,-0.03125,-0.0078125,-0.03125,0.015625,-0.0546875,-0.0078125,0.078125,0.0234375,-0.0234375,0.0234375,-0.0078125,0.0625,0.0390625,-0.03125,0.03125,-0.015625,-0.0625,0.015625,-0.0546875,-0.0390625,0.1015625,0.0390625,-0.0546875,0.046875,0.0390625,0.0078125,0.0078125,0.015625,-0.0078125,-0.0078125,-0.03125,-0.078125,-0.0390625,-0.0078125,-0.046875,0.015625,0,0.0078125,-0.0703125,0.0546875,-0.0078125,0.0546875,-0.015625,0.0390625,0,0.0078125,-0.0078125,0,0.015625,0,0,0,0,-0.015625,-0.0390625,0.046875,0.0078125,-0.046875,0.0546875,-0.0234375,-0.1328125,-0.0703125,-0.0078125,-0.0234375,0,0.0625,-0.03125,0.0625,-0.078125,-0.0078125,-0.0390625,0.0390625,0.0546875,0.03125,-0.09375,-0.0390625,-0.03125,0.015625,0.046875,0.140625,0.0078125,0.015625,0,0,0,0,-0.0078125,-0.015625,0,-0.03125,0.0546875,0.03125,-0.015625,-0.0234375,0.0625,0.0703125,-0.015625,-0.0625,-0.03125,0.0078125,-0.015625,0.0234375,-0.046875,-0.015625,0.046875,-0.046875,0.0546875,0.0078125,-0.0625,-0.03125,-0.0078125,-0.0703125,-0.0078125,-0.0078125,-0.015625,0.015625,0.0078125,-0.03125,0,-0.0078125,0.0234375,0,0.0390625,-0.109375,-0.03125,-0.0078125,-0.0078125,-0.0859375,0.046875,0.0625,-0.0390625,-0.078125,-0.0703125,-0.0390625,-0.0078125,0.0078125,0,-0.0390625,0.0078125,0.0078125,0.0546875,0.03125,-0.015625,-0.0390625,0.015625,0.0078125,0.0078125,-0.0390625,0.03125,0.0078125,-0.0546875,-0.015625,0.0234375,0.0078125,0,-0.0078125,-0.0390625,0.0546875,0.015625,0.0625,0.015625,-0.0234375,0.015625,-0.0078125,0.0078125,-0.0234375,-0.03125,0.0859375,-0.0390625,0.0703125,0.03125,0.0390625,0.0390625,-0.0234375,-0.0859375,-0.078125,0.046875,-0.0546875,0.015625,0,-0.0078125,-0.0078125,0,0.0078125,0.0078125,0,-0.015625,0.0078125,0,-0.0078125,0.0234375,0.03125,0,0.0078125,0,-0.046875,0.0078125,-0.0546875,-0.015625,-0.046875,0.0078125,-0.0546875,0.1015625,-0.1328125,-0.015625,0.0234375,0,0.015625,0.0078125,-0.015625,-0.0234375,0.03125,0.109375,0.046875,-0.0234375,-0.015625,0.0234375,-0.0078125,-0.0546875,-0.0234375,0.0078125,-0.0546875,0.0390625,0.0390625,0,-0.0078125,-0.0390625,-0.1015625,-0.046875,-0.0078125,0.1015625,-0.015625,-0.0078125,0.0625,-0.0390625,0,-0.0625,0.0234375,-0.015625,0,0.046875,-0.0703125,-0.015625,-0.0546875,-0.0546875,0,0.03125,0.0234375,-0.15625,0.078125,-0.03125,0.0546875,0.015625,-0.03125,-0.0234375,0.0546875,-0.0546875,-0.0703125,0.0234375,-0.0625,0.0390625,-0.0234375,0.0078125,0.046875,-0.0078125,-0.1015625,0.015625,0.015625,0,0.03125,0.03125,0.0078125,0.0390625,-0.09375,0.0390625,0.046875,-0.0546875,-0.015625,-0.015625,-0.0390625,-0.03125,0.0390625,-0.1484375,0.0546875,0.0546875,-0.0703125,0.078125,-0.046875,0.0078125,-0.046875,-0.0390625,0.0703125,0.109375,-0.0234375,-0.0234375,0.09375,-0.0234375,-0.0390625,-0.03125,0.125,-0.03125,0.03125,-0.0390625,-0.015625,-0.125,-0.0390625,-0.0078125,-0.015625,0.046875,0.1015625,-0.0390625,-0.0546875,0.0546875,-0.0625,-0.015625,0,0.0390625,0.0078125,0.0625,-0.03125,-0.0234375,0.0078125,-0.0234375,0.0234375,-0.015625,-0.0078125,0,0.078125,-0.0234375,-0.0234375,0.078125,0.03125,0,-0.0078125,-0.015625,0.0078125,-0.0078125,0.0078125,-0.0078125,0.0078125,0.015625,0.0078125,-0.0234375,0.0078125,0.015625,-0.0546875,-0.0625,0.0234375,-0.0234375,0.0859375,0,-0.0234375,0.015625,0.0078125,0.03125,-0.0078125,-0.03125,-0.0078125,-0.0234375,-0.015625,0.0078125,-0.015625,-0.0078125,-0.0234375,-0.015625,-0.0078125,-0.0078125,0.0703125,0.0078125,0,0,0,0,0,0.0078125,0.0078125,-0.015625,-0.0234375,-0.03125,-0.0078125,-0.0234375,0.03125,0.0234375,0,-0.0078125,-0.0078125,0,0,-0.046875,-0.0234375,-0.046875,0.0390625,-0.0390625,0.0234375,0.09375,0,0.046875,0.0234375,-0.0078125,-0.0234375,-0.046875,-0.0234375,-0.1015625,0.0390625,0.015625,-0.03125,-0.0234375,-0.0078125,-0.0625,-0.0390625,-0.0078125,0,0.015625,0.0078125,-0.0234375,-0.0234375,-0.0234375,0.03125,0.046875,-0.0078125,-0.0078125,0,0,0,-0.0234375,-0.03125,0.0078125,0,0,0.0234375,0.0625,0.015625,0.0078125,0,0.015625,0,0.0234375,0.0078125,0.0078125,0.0078125,0.0078125,0.0078125,0.0078125,0.0078125,-0.0078125,-0.015625,0.0390625,-0.0390625,-0.0546875,0,0.015625,-0.0234375,-0.015625,0.0078125,0.0078125,-0.015625,0.0859375,-0.0390625,-0.015625,-0.015625,-0.0078125,-0.0234375,-0.0390625,0.0078125,0.0390625,-0.015625,-0.03125,-0.0078125,0,0,0.0078125,-0.0078125,0.0078125,0.0078125,0.0078125,0.0234375,0.015625,-0.0078125,-0.0234375,-0.015625,-0.015625,-0.0078125,0.0078125,-0.0390625,0.0078125,-0.015625,-0.015625,0.0234375,-0.015625,-0.0234375,-0.0546875,0,-0.0078125,-0.0234375,-0.0078125,-0.0390625,-0.03125,-0.03125,-0.0234375,0.0234375,-0.0234375,-0.0234375,0.078125,0,-0.0078125,-0.015625,-0.0390625,-0.0859375,-0.046875,0.0234375,0.0078125,-0.046875,0.015625,-0.015625,-0.0390625,-0.015625,0.03125,0,0.03125,0.03125,0.03125,0,0.0234375,0.015625,0.015625,-0.0234375,-0.03125,0.0234375,0.03125,0.0390625,-0.015625,-0.0078125,-0.0234375,-0.015625,-0.0546875,0,0,-0.0703125,0.0625,0.0078125,-0.0078125,0.015625,-0.0078125,-0.046875,-0.03125,-0.015625,-0.015625,0.0078125,-0.015625,0.015625,0,0.0078125,0.0234375,-0.0234375,-0.0078125,0,0,0,-0.03125,-0.0234375,-0.0234375,0,0.1015625,0.0390625,-0.03125,0.015625,-0.015625,0.015625,-0.0234375,-0.0234375,0.015625,-0.0625,0.015625,0.0546875,-0.0703125,0.0078125,0,-0.0078125,-0.0078125,-0.0078125,-0.015625,-0.03125,-0.0234375,-0.03125,-0.015625,0,0,0.015625,-0.015625,0.03125,0.015625,0,-0.0625,-0.015625,0,-0.015625,0.03125,-0.03125,0.0078125,0,-0.046875,0,0.0078125,-0.0078125,-0.03125,-0.046875,0.046875,0,-0.0078125,-0.015625,0.0390625,-0.0078125,-0.046875,-0.0703125,0.0390625,-0.046875,0.046875,0.1015625,0.0234375,-0.0078125,-0.0078125,-0.0078125,0.0078125,-0.015625,-0.0078125,-0.0234375,0.0078125,0,-0.0078125,0.03125,0,-0.03125,-0.09375,-0.1015625,0.015625,-0.0078125,-0.03125,-0.0078125,0.015625,-0.015625,-0.0703125,0.0078125,-0.0390625,-0.0390625,-0.0078125,-0.046875,0.0078125,-0.046875,0.0078125,0.0546875,-0.0078125,-0.0078125,-0.046875,-0.0234375,0.09375,-0.125,-0.0078125,-0.015625,0.0078125,0.0078125,0.0078125,0.015625,0.0078125,0,0.0078125,-0.0546875,-0.0390625,0.015625,0.0078125,-0.03125,-0.0390625,0.03125,0.0859375,-0.078125,0.1484375,0.078125,-0.046875,0.046875,-0.0625,-0.0390625,0.0625,-0.015625,-0.015625,-0.0234375,-0.0078125,-0.09375,-0.0078125,-0.0546875,-0.0078125,0.078125,0.078125,-0.0703125,-0.0078125,0.0078125,0,-0.0078125,-0.0078125,0.0078125,-0.0390625,0.0078125,0.0078125,-0.0390625,0.0078125,0.015625,0.015625,0.03125,0.1015625,-0.046875,-0.0390625,-0.0078125,-0.03125,-0.0625,0.0390625,0.0625,0.0625,-0.0234375,0,-0.0625,0.015625,-0.0234375,0.09375,-0.015625,-0.0234375,0,0,-0.046875,0.0078125,0.0078125,-0.046875,-0.0234375,-0.046875,0.0546875,0.0234375,-0.0390625,-0.046875,0.0234375,0.015625,-0.015625,0.015625,0.0390625,0.078125,0.015625,0.046875,-0.0390625,-0.0390625,-0.0234375,0.0546875,-0.0703125,0.109375,0.0078125,-0.140625,-0.0078125,0.0390625,0.0546875,-0.0234375,-0.0078125,-0.015625,-0.03125,-0.015625,-0.0234375,-0.0234375,0.0078125,0,-0.0078125,-0.0078125,-0.0078125,-0.0390625,0.015625,0.0703125,-0.046875,-0.0546875,-0.0078125,0.0546875,0.03125,-0.015625,-0.0625,-0.0859375,-0.0078125,-0.0078125,0,-0.0234375,0.046875,-0.015625,-0.015625,0.0390625,-0.0234375,-0.03125,-0.0546875,0.0625,0.125,-0.0625,-0.0078125,0.0078125,0.046875,-0.1171875,-0.046875,-0.015625,-0.046875,-0.0546875,0.0546875,-0.0625,-0.0546875,-0.0390625,-0.0390625,-0.0234375,0.0078125,0.0390625,-0.0390625,-0.0234375,0.0625,-0.0703125,0.03125,-0.0625,-0.0078125,0.0546875,0.0234375,0.0390625,0,0.078125,0,0.0078125,-0.0234375,-0.0078125,0.0390625,-0.078125,-0.078125,0.140625,-0.09375,-0.0703125,0.0703125,-0.0546875,0.0546875,0.0703125,-0.1015625,-0.0703125,0.046875,0.0390625,0.0078125,0.046875,-0.015625,-0.0234375,0.0625,0.0234375,0.0390625,0,-0.0859375,-0.0390625,-0.0078125,0,0.03125,0,0,0.1328125,-0.015625,0.0859375,0.03125,0.015625,-0.0078125,-0.015625,-0.0390625,-0.015625,-0.0390625,0,-0.0234375,-0.09375,0.0546875,0.015625,-0.0078125,-0.109375,-0.0390625,-0.1171875,-0.015625,0.0703125,0.1328125,-0.0546875,-0.03125,0.0546875,-0.1015625,-0.078125,0.03125,0.03125,0.0625,-0.0390625,0.125,0.0078125,-0.03125,-0.015625,0.0078125,0.015625,0.0234375,0.046875,0.015625,-0.0390625,0.0078125,-0.1640625,-0.0625,-0.0234375,-0.046875,-0.0234375,-0.015625,-0.03125,-0.0546875,-0.078125,-0.015625,0,0.078125,0.0703125,0.0390625,-0.0078125,-0.015625,0.015625,-0.0078125,0.0078125,0,0.015625,-0.0078125,0,0.0078125,-0.0234375,-0.03125,-0.0078125,-0.078125,0.0703125,0.0625,-0.0390625,-0.0390625,0.0625,0.0390625,-0.0859375,-0.0234375,-0.0390625,-0.0546875,0.015625,0.03125,-0.0390625,0,-0.015625,0.046875,0.03125,-0.03125,0.078125,-0.03125,-0.0390625,0.0078125,-0.0078125,0.0078125,0.0078125,-0.0078125,0,0.0078125,0.015625,0.0078125,-0.0078125,0.0078125,-0.0234375,0.0234375,-0.0078125,0.0078125,0.015625,0.0234375,0,0,0.0390625,-0.1640625,-0.015625,0.0078125,-0.0078125,-0.0625,-0.0078125,0.0234375,0.015625,-0.046875,-0.03125,-0.0234375,0,-0.0703125,0.0546875,-0.0234375,-0.0234375,-0.0234375,-0.0390625,-0.0078125,0.1171875,0.0078125,-0.015625,0,0.0234375,-0.0234375,0.0078125,0.015625,0,-0.0234375,-0.0390625,0.015625,-0.0703125,-0.03125,-0.0625,-0.03125,-0.03125,-0.015625,-0.0078125,0.046875,0.03125,-0.015625,0.0078125,-0.0234375,-0.0234375,0,0.0234375,-0.03125,-0.015625,-0.0546875,0.0078125,0.0234375,-0.0078125,0,-0.0234375,0.0234375,-0.0234375,0.0703125,-0.0625,-0.0078125,0.0234375,-0.0234375,-0.0234375,-0.03125,0.03125,0.0234375,0.0234375,-0.0078125,-0.0234375,-0.03125,0.0078125,-0.0390625,0.03125,0.109375,0.0390625,-0.03125,-0.046875,0.0546875,0.015625,-0.0859375,-0.0078125,0,0.015625,0.0078125,-0.0234375,0.0234375,0,0.0078125,0.015625,-0.0234375,-0.0234375,-0.0625,-0.03125,-0.0078125,-0.0078125,0.0078125,-0.0078125,0.03125,0,0.0546875,-0.015625,0,0.078125,-0.03125,0,0,0.015625,-0.0078125,-0.0078125,-0.0703125,0.046875,0.0234375,-0.09375,-0.0234375,-0.015625,-0.0625,-0.0625,0.0078125,-0.1171875,0.0546875,0.0625,0.0859375,0.03125,-0.03125,-0.015625,-0.03125,-0.0546875,-0.046875,0.0390625,-0.0234375,-0.03125,0.0078125,-0.0390625,0,-0.0234375,-0.0390625,0.0859375,-0.0703125,-0.015625,-0.0234375,0.0703125,-0.015625,0.015625,-0.0234375,0.0703125,0.1640625,-0.078125,-0.046875,-0.0390625,0,0,0.0234375,-0.0546875,0.015625,-0.0546875,-0.0546875,0,0,0.015625,0.0078125,-0.0078125,-0.0078125,-0.015625,0.0078125,-0.03125,0.015625,-0.0625,-0.0078125,-0.0703125,-0.015625,0.0078125,-0.0078125,-0.0546875,-0.03125,0.046875,0.0703125,0,0.0078125,-0.0703125,-0.015625,-0.1484375,-0.0234375,-0.09375,-0.0234375,0.0390625,0.015625,0.0546875,-0.0625,0,0,-0.0390625,0.0625,0.0234375,0.0234375,-0.0078125,-0.0234375,-0.0625,0.015625,0.0625,0.1171875,-0.015625,0.0234375,-0.015625,-0.0390625,-0.0234375,-0.0078125,-0.015625,-0.1015625,0.0234375,0.0078125,0.015625,0.0390625,0.0546875,0.03125,0.0078125,0.0234375,0.0078125,0.0078125,-0.09375,-0.03125,-0.0859375,-0.046875,0.0078125,0.0859375,0.015625,0.015625,0.0625,0.03125,0.09375,-0.03125,0.015625,0.0390625,-0.015625,-0.0234375,-0.015625,-0.015625,0.0078125,0.015625,0.0078125,-0.0078125,0.015625,0.0078125,-0.015625,-0.0390625,-0.015625,0.1328125,-0.03125,-0.0078125,-0.0234375,0.0703125,0.015625,-0.0078125,-0.0078125,0.015625,0,0.03125,0.0234375,-0.03125,0.03125,-0.0234375,0.0078125,-0.0625,-0.015625,-0.0234375,-0.0390625,-0.0390625,-0.03125,0.03125,-0.015625,-0.0234375,-0.0078125,-0.0078125,-0.015625,-0.015625,0.0078125,0.0078125,0,-0.015625,0.0078125,-0.0546875,-0.0625,-0.015625,-0.0078125,0.0390625,-0.015625,-0.109375,-0.0078125,-0.0234375,-0.125,0.0859375,-0.0390625,0.046875,-0.0703125,-0.03125,0.1484375,0.0234375,-0.0390625,-0.0859375,-0.0234375,-0.015625,0.03125,-0.015625,-0.0078125,0.1015625,-0.078125,-0.0390625,0.0390625,0.1015625,0.0078125,-0.03125,0,-0.0078125,-0.046875,-0.015625,0.0234375,-0.0703125,-0.046875,-0.03125,-0.0234375,0.0390625,-0.0234375,-0.046875,-0.0625,-0.03125,-0.046875,0.0078125,0,0,0,-0.0390625,0.09375,-0.09375,-0.0078125,-0.03125,0.0234375,0,-0.0390625,-0.015625,0.015625,0.0078125,0.0078125,-0.015625,0.03125,-0.0234375,-0.015625,0.0390625,-0.0390625,0.015625,-0.015625,-0.015625,-0.015625,0.0625,0.171875,0,-0.125,-0.0859375,-0.046875,-0.03125,0,-0.0390625,-0.0625,0.0078125,-0.046875,0.0625,0.0234375,0,-0.0234375,-0.0234375,-0.015625,0.0078125,0.0078125,-0.0078125,0,-0.03125,-0.0078125,0.015625,0.0078125,0,-0.015625,-0.015625,0.0234375,-0.046875,-0.0390625,0.0234375,0.0546875,0.0078125,0,0.0546875,-0.0390625,0,0.0234375,-0.0078125,-0.0390625,0.0234375,0.0078125,-0.0234375,-0.0078125,0.046875,-0.0390625,-0.078125,-0.0234375,-0.03125,0.1484375,-0.0234375,-0.0234375,0.0625,-0.09375,-0.0390625,-0.078125,0.09375,-0.0078125,-0.03125,-0.0390625,0.0078125,-0.09375,0,0.0234375,-0.1171875,0.046875,0.046875,0.0859375,-0.0234375,-0.0546875,0.015625,-0.046875,0.0234375,0.0546875,-0.09375,-0.03125,0.0703125,-0.015625,-0.0546875,0.0703125,0,0.03125,-0.0078125,-0.125,-0.0078125,-0.015625,-0.046875,-0.0703125,-0.0625,-0.015625,-0.0078125,-0.1015625,0.046875,-0.0078125,0.1015625,0.0234375,0.015625,0,-0.015625,0,-0.0078125,-0.0546875,-0.015625,0.1171875,-0.0078125,-0.0234375,-0.0859375,0.03125,0.046875,0.0390625,-0.0390625,-0.0390625,0.03125,-0.078125,-0.046875,0.0390625,0,-0.03125,0.0625,0.046875,-0.0078125,-0.0234375,-0.0625,-0.0390625,-0.0546875,0.0078125,0.0859375,-0.0625,0.0625,-0.0625,-0.0234375,-0.015625,0.0078125,-0.03125,0.0234375,0.03125,0.0234375,-0.171875,-0.0234375,-0.03125,0.1328125,-0.046875,-0.015625,-0.078125,-0.0625,0.0703125,-0.0703125,-0.0390625,0.03125,0.0234375,-0.03125,0.015625,0,0.0546875,0,-0.0703125,0.0078125,0.0390625,-0.046875,-0.046875,-0.0078125,0.046875,-0.0546875,-0.0859375,-0.0625,0.015625,0.0234375,-0.03125,-0.03125,-0.015625,-0.015625,0.015625,0.0078125,-0.0078125,-0.0078125,0.0234375,0,0,0,0.015625,-0.0390625,0.0078125,0,-0.0078125,0.0234375,-0.03125,0.015625,-0.0078125,0.015625,-0.015625,-0.0078125,0.03125,-0.0078125,0,-0.046875,-0.03125,0.0078125,-0.0546875,-0.0234375,-0.0546875,-0.03125,0.0390625,-0.0078125,0.0546875,-0.0546875,0,0,0.0078125,0.015625,-0.0078125,0.0078125,0,0.0078125,-0.0078125,-0.0625,0,-0.0078125,-0.09375,0.03125,0.0234375,0.015625,-0.0390625,-0.078125,0.0703125,0.0703125,0.046875,0.0234375,-0.015625,0.078125,-0.0390625,-0.03125,-0.0390625,0.0625,0.0625,-0.0546875,-0.0546875,-0.015625,0.0078125,-0.03125,-0.0390625,-0.046875,-0.03125,0.0390625,0.03125,-0.0390625,0.0078125,0.0625,-0.015625,-0.015625,-0.015625,-0.0234375,0.0078125,-0.0234375,0,-0.0625,0.0390625,-0.0234375,-0.03125,-0.0390625,-0.0078125,-0.0546875,0.0390625,-0.0234375,0.0390625,-0.0078125,0.03125,0.0234375,0,0.03125,0.0390625,-0.0078125,-0.0078125,0.0078125,0.0390625,-0.0234375,-0.015625,0,0.03125,0.0078125,-0.0234375,-0.03125,-0.0546875,-0.0234375,0.0234375,-0.0078125,0.0078125,-0.03125,-0.09375,0,-0.0234375,-0.015625,0.0234375,0.0625,-0.0234375,-0.0625,0.015625,0,0.078125,0.0078125,0,-0.046875,0.015625,-0.0859375,-0.03125,0,-0.0078125,-0.015625,-0.0078125,-0.0078125,-0.03125,0,0.0078125,0,-0.0078125,-0.0546875,-0.03125,0.0390625,0.046875,-0.03125,0.015625,-0.03125,-0.015625,-0.0234375,0.0234375,0.0234375,0,0.0078125,0.015625,-0.015625,0,0.0078125,0.03125,0,0.0859375,-0.0390625,-0.0234375,0.0625,-0.0234375,-0.015625,-0.0390625,0,-0.0390625,0.046875,-0.078125,0.0078125,0.0078125,0.03125,0,-0.0234375,0.0234375,0,0.015625,-0.0390625,-0.0546875,-0.015625,-0.0390625,-0.0234375,-0.03125,0.0078125,0.0234375,-0.0390625,0.0390625,0.0625,0.0390625,-0.0390625,-0.015625,-0.0078125,0.046875,0.0234375,-0.015625,0.0859375,-0.046875,-0.0078125,-0.03125,0.015625,0,0.03125,-0.0625,0.015625,0.0625,0.015625,-0.0234375,0.03125,-0.0234375,-0.015625,0.0703125,0,-0.0234375,0.09375,-0.046875,-0.0078125,-0.03125,-0.0234375,0.015625,-0.0390625,0.0078125,0,-0.03125,-0.0625,-0.046875,-0.03125,-0.0078125,-0.0078125,-0.0859375,-0.03125,-0.0703125,-0.0234375,0,-0.015625,0.0859375,0.03125,0.0078125,-0.0390625,0.078125,-0.0390625,0.0078125,-0.0078125,0.0625,-0.0234375,-0.0234375,-0.015625,-0.0390625,0.046875,-0.03125,0.03125,-0.0625,-0.0390625,-0.015625,-0.0390625,-0.015625,-0.0390625,0.0078125,0.0078125,0,-0.0234375,0.0625,-0.015625,-0.0078125,0.046875,0,0.0078125,0,0.0625,-0.078125,0.0625,-0.015625,-0.0234375,-0.03125,0,0.0234375,0.0078125,-0.03125,0.0390625,0.0390625,-0.0625,0.0390625,0.0234375,-0.0078125,-0.0078125,-0.0078125,-0.0078125,-0.015625,-0.0078125,0,0.015625,-0.0078125,-0.03125,-0.0234375,0.0625,-0.0234375,-0.0703125,0.0078125,-0.0078125,0,0.0078125,-0.0234375,-0.015625,0.0078125,0,-0.015625,0.046875,0.0234375,-0.0078125,0.0078125,0.109375,0.1015625,-0.0546875,-0.0234375,-0.0625,-0.015625,-0.0234375,-0.09375,0.015625,0.0078125,-0.0078125,-0.0078125,0,0.0078125,0.0078125,0,0.0078125,-0.015625,0.0390625,-0.0234375,0.0546875,0.0234375,-0.0234375,0.0234375,-0.0234375,0.015625,0,0,0.078125,-0.015625,-0.0234375,-0.0625,-0.0625,-0.0078125,-0.015625,0.015625,0.09375,0.1171875,-0.03125,-0.109375,-0.0078125,-0.0078125,-0.0234375,-0.03125,0.015625,-0.0546875,-0.03125,0,-0.0234375,-0.0234375,-0.015625,0.0390625,0.0390625,-0.015625,-0.0234375,-0.03125,0,-0.0546875,-0.03125,-0.0078125,-0.0234375,-0.015625,-0.03125,0.015625,-0.0078125,-0.03125,0.015625,0,0.0234375,-0.0234375,0.0078125,0.015625,0.0546875,0,-0.0546875,0.015625,0.03125,-0.0078125,0,0,0.0234375,0.03125,0.0234375,-0.0078125,-0.046875,0,0.0078125,0.0234375,0.0078125,0.0234375,-0.015625,0.03125,-0.046875,0,-0.0703125,-0.0078125,-0.0234375,0.0234375,-0.0078125,-0.03125,0.046875,-0.015625,-0.0078125,0.015625,-0.0078125,-0.0078125,0.015625,-0.03125,-0.015625,0,0,0,0.0078125,0.0078125,0,0.015625,0.015625,0.0078125,-0.03125,0.0078125,0.0234375,0,-0.015625,-0.015625,0,0,0.0078125,0.046875,0.0546875,-0.015625,-0.0078125,-0.0546875,-0.0234375,-0.015625,-0.03125,-0.015625,0.0625,-0.0234375,-0.03125,-0.046875,0.015625,0.015625,0.03125,-0.015625,0.046875,0.078125,0,-0.015625,-0.0625,-0.0625,0.0078125,-0.0078125,0.015625,-0.015625,-0.0859375,-0.1015625,0.015625,-0.015625,-0.03125,-0.0234375,0.0546875,-0.015625,0,-0.0546875,-0.03125,-0.015625,-0.015625,0,-0.0390625,-0.03125,0.0078125,0.0625,0.0078125,-0.0390625,0.015625,-0.1015625,-0.0078125,0.0546875,0.0078125,0.0078125,-0.0234375,0.0078125,-0.015625,0.0703125,-0.046875,-0.0625,-0.03125,-0.046875,-0.015625,0.0859375,0.046875,-0.0390625,0.03125,-0.078125,-0.015625,-0.046875,-0.046875,0.0234375,0.0078125,0.0546875,-0.0078125,-0.0234375,0.03125,0,-0.0546875,0.0078125,0.0703125,0.140625,0.0078125,-0.015625,0.0078125,0.046875,0,-0.0390625,-0.03125,0.0234375,0.046875,-0.0859375,0.0546875,-0.046875,-0.0078125,-0.0625,0.015625,0.03125,-0.015625,-0.03125,-0.046875,-0.0078125,-0.015625,0.09375,-0.0234375,-0.015625,0.015625,-0.046875,-0.0234375,-0.015625,-0.015625,-0.015625,-0.0078125,-0.0078125,0.0234375,-0.0234375,-0.0390625,0.0078125,-0.03125,-0.0546875,-0.03125,0.0546875,-0.046875,-0.0390625,0,0,0,-0.0078125,0.0078125,-0.0234375,0.015625,0.03125,-0.0078125,-0.0078125,-0.078125,0.0078125,0,-0.0078125,-0.0078125,0.0078125,0.0078125,0,-0.0078125,0.015625,-0.0078125,-0.0546875,0,-0.0234375,-0.0390625,0.0390625,-0.015625,-0.0546875,0.015625,0.0078125,0.0078125,0,0.0078125,-0.0078125,0.0078125,-0.015625,-0.0390625,-0.0390625,0,0,0.03125,-0.015625,-0.0078125,0.03125,-0.015625,0.0234375,0.0078125,0.0078125,0,-0.015625,0.015625,-0.0078125,0.0078125,0,0.015625,-0.0078125,0.0078125,-0.015625,0,0,-0.0078125,-0.0234375,-0.0234375,0.0625,-0.015625,-0.0234375,0.015625,0.046875,-0.0234375,-0.0390625,0.0390625,0,0.0234375,-0.0859375,-0.0234375,0.0234375,-0.0234375,-0.015625,-0.0546875,-0.03125,-0.0234375,-0.03125,0.015625,-0.0078125,-0.0390625,-0.015625,0,-0.0390625,0.0703125,-0.015625,0,-0.0234375,0.015625,0.015625,0.03125,-0.0078125,-0.0390625,-0.0390625,0,0.046875,0,0.015625,-0.0390625,0.015625,-0.015625,0.0390625,0.015625,-0.0078125,0.0078125,-0.046875,0.0078125,0,0.0390625,0,-0.0078125,-0.015625,0,0.015625,0,-0.0078125,0,0,-0.015625,-0.015625,0.015625,-0.0234375,0.0078125,0.015625,-0.0078125,-0.046875,-0.03125,-0.0234375,-0.0234375,-0.0078125,0.0078125,0.0625,0.03125,0,0,-0.0234375,-0.015625,0.0078125,-0.0390625,-0.0078125,0.0234375,0.0390625,0.0078125,0.0078125,0,-0.0078125,0.015625,0.0078125,0,-0.0078125,0.0234375,0,-0.03125,0,-0.015625,-0.0078125,0,0,0,0.03125,0.0078125,0,-0.0078125,0,-0.0078125,-0.046875,-0.0078125,0.0703125,0.0078125,-0.015625,-0.0390625,-0.0625,0.015625,-0.0390625,0.046875,-0.0078125,0,0.015625,-0.0078125,0.015625,0,-0.0078125,-0.0390625,-0.109375,-0.0234375,0.03125,0.046875,-0.0078125,0.0390625,0.0234375,-0.015625,0,-0.078125,-0.03125,0.015625,0.046875,0.0078125,0.0078125,0,0,0.015625,0.015625,-0.0234375,-0.0546875,0,-0.015625,-0.015625,-0.046875,-0.015625,0.015625,0.0625,0,-0.09375,-0.015625,-0.0078125,-0.03125,-0.0390625,-0.0078125,-0.0078125,0.03125,0.0078125,-0.015625,0.046875,-0.0078125,0.0390625,0.0234375,-0.0078125,-0.0234375,-0.046875,0,-0.0703125,-0.015625,0,-0.0703125,0.078125,0,-0.0078125,-0.046875,-0.0234375,0.03125,-0.0234375,-0.015625,-0.0078125,-0.0546875,-0.03125,0.0390625,-0.09375,-0.015625,0,0.0390625,-0.015625,-0.0078125,0.015625,0,0.015625,0,-0.0078125,0.0625,0.0390625,-0.0078125,-0.046875,0.0234375,-0.015625,0.0234375,0.0078125,-0.0078125,-0.03125,-0.0625,0,-0.0078125,0.046875,-0.015625,0.0625,0.0703125,-0.0234375,-0.015625,0.0234375,0.0078125,0.0546875,0.0390625,-0.015625,0.0234375,0,-0.015625,-0.0390625,-0.015625,-0.0234375,0.0234375,-0.0234375,-0.03125,0.0625,0.0234375,0.0625,0.0234375,-0.0078125,-0.0078125,0,0,0.0078125,-0.0078125,-0.0078125,-0.0078125,-0.0078125,0,0.046875,0.03125,-0.0234375,0.015625,-0.015625,0,0.0234375,0.0390625,-0.015625,0.0078125,-0.0390625,-0.0546875,0.0234375,-0.1015625,0.0234375,-0.0625,0.046875,-0.03125,0.0703125,0.0703125,-0.015625,0.03125,-0.0390625,0.0234375,0.0703125,-0.0390625,-0.03125,0,0.0078125,0,0.015625,-0.0078125,0.0078125,-0.0078125,-0.0078125,0,-0.015625,0.046875,-0.03125,0,-0.0859375,-0.03125,-0.0078125,-0.0859375,-0.03125,0.0546875,0,0,-0.0234375,0.0390625,-0.0078125,0.0234375,0.0078125,-0.0234375,0.0234375,0.046875,-0.0234375,0.015625,0,0.0234375,0.0078125,-0.046875,-0.0390625,-0.046875,0.0546875,0.015625,-0.015625,0.015625,0.0078125,-0.015625,-0.0234375,-0.0078125,0.0703125,0.03125,-0.0703125,-0.03125,0.0078125,-0.0234375,0,0.0234375,-0.0234375,-0.015625,0,0.0390625,0.0390625,-0.015625,-0.0078125,0,-0.03125,0,0.0234375,-0.0078125,-0.015625,0,0.0078125,-0.0234375,0,-0.015625,0,0,-0.015625,0.0625,-0.0390625,-0.0625,-0.0078125,-0.0390625,0.015625,-0.015625,0.0078125,0.046875,-0.03125,-0.0078125,0.0078125,-0.0390625,-0.015625,-0.03125,0,0.0234375,0.0078125,0.015625,0.0625,-0.0078125,-0.015625,-0.015625,-0.0859375,-0.015625,0.015625,-0.0078125,-0.0078125,-0.015625,0.015625,0.0078125,0.0078125,0,-0.015625,-0.0078125,-0.0703125,-0.0078125,-0.0625,-0.03125,-0.0234375,0.0078125,-0.015625,-0.0078125,-0.0078125,-0.0390625,0.0078125,-0.0546875,0.046875,-0.015625,-0.0546875,0.0546875,-0.0390625,0,0.0546875,0,0.0625,-0.0234375,0.0390625,-0.03125,-0.0546875,0.0078125,-0.03125,0.0078125,-0.0390625,-0.015625,-0.0234375,-0.0390625,-0.046875,-0.0078125,-0.015625,0.046875,-0.0546875,-0.0390625,-0.1015625,-0.0078125,0,-0.0625,-0.0234375,-0.0234375,0,0.015625,-0.015625,0.015625,0.046875,-0.0234375,0.046875,0.046875,-0.015625,-0.0546875,-0.078125,0.0546875,0.0546875,-0.015625,0,0.03125,0,-0.0390625,-0.0078125,-0.0546875,-0.0078125,-0.0078125,-0.0234375,-0.0234375,0.0625,-0.0625,0,-0.03125,-0.015625,-0.0078125,-0.0390625,-0.015625,-0.03125,0.171875,-0.0234375,-0.0078125,-0.015625,0.0078125,0,0.0390625,-0.0625,0.0859375,0.0234375,0.0234375,-0.03125,-0.0390625,-0.0625,0.1015625,-0.0703125,0.03125,-0.0546875,0,0.0234375,-0.03125,-0.0546875,-0.03125,-0.015625,0,-0.078125,-0.0390625,-0.0703125,-0.0703125,-0.015625,-0.0078125,0.0078125,-0.0390625,-0.046875,-0.0546875,-0.0078125,-0.0703125,0.0390625,-0.0234375,0,-0.0078125,-0.015625,0.046875,0.0859375,-0.0078125,-0.015625,-0.015625,0,-0.1171875,0.015625,-0.03125,-0.0625,-0.0546875,-0.0078125,0,0.046875,-0.015625,0.0390625,0.0078125,0.078125,-0.03125,-0.015625,-0.0078125,0.03125,0,0.0703125,-0.0078125,-0.0078125,-0.0078125,0.015625,0,0.0078125,-0.0078125,0.015625,-0.0078125,0.015625,-0.0078125,-0.1328125,-0.03125,-0.015625,-0.1015625,0.0390625,-0.0078125,0.0234375,0.0078125,0.0234375,-0.015625,-0.015625,0.046875,-0.0859375,0.0546875,0.0234375,0,-0.0234375,0.0078125,0.03125,-0.0078125,-0.078125,0,-0.0390625,-0.0390625,-0.0390625,0,-0.015625,-0.0078125,0,0.015625,0,0,-0.0078125,-0.0078125,-0.03125,-0.0234375,-0.046875,-0.046875,0.03125,-0.0234375,-0.03125,-0.03125,-0.0078125,0.078125,0.0390625,-0.0234375,0.0390625,-0.0390625,-0.0703125,-0.015625,0.0390625,0.0625,-0.0234375,-0.0703125,-0.0390625,0,-0.0234375,0.03125,-0.0234375,-0.03125,0.046875,0,0.0234375,-0.015625,-0.0078125,-0.0234375,0.0234375,0.0234375,0,0.0234375,-0.0078125,-0.015625,0.0703125,0.0078125,-0.03125,-0.03125,-0.015625,0.0390625,0.03125,0,0,0,-0.015625,-0.015625,-0.046875,-0.03125,0.015625,0.0390625,-0.015625,-0.0390625,-0.0078125,0,-0.0078125,-0.03125,-0.015625,0.0390625,0.0234375,-0.0078125,-0.078125,-0.0078125,0.0234375,-0.0078125,0.0234375,0,-0.03125,-0.0703125,0,0.1015625,0.1015625,0,-0.0078125,-0.0703125,0,0.0703125,-0.0234375,-0.015625,-0.0234375,-0.0078125,0.0234375,-0.0078125,0.125,0.0078125,-0.015625,-0.046875,0,-0.015625,-0.0078125,0,0.0078125,0.015625,0,0.0078125,-0.015625,-0.0078125,0,-0.0234375,-0.015625,0.015625,0,-0.015625,-0.0234375,0.046875,0.03125,0.0546875,0.015625,0.015625,0.03125,0,-0.0234375,0.1015625,-0.015625,0.0078125,0.015625,0.109375,0.015625,-0.0703125,-0.046875,0,0,0.0703125,-0.0078125,0.0234375,0.1015625,-0.0234375,0.0390625,-0.0390625,-0.0234375,0.015625,-0.046875,-0.0078125,0.015625,0.015625,-0.0078125,-0.0078125,0.03125,-0.0390625,-0.03125,0.09375,0.0234375,-0.0234375,-0.0234375,-0.0546875,0,0.0078125,-0.0078125,0.015625,-0.0234375,0.015625,0.0546875,0,0.015625,-0.0078125,-0.0625,0.0390625,0.0234375,-0.0234375,-0.03125,-0.0390625,0.046875,-0.015625,-0.0234375,0.09375,-0.015625,0.03125,0.0234375,0.0234375,0.0234375,0.015625,0,-0.046875,-0.0078125,0,-0.0703125,-0.0703125,0.0234375,-0.0234375,0.0390625,-0.0078125,0.0390625,0.03125,-0.015625,0.015625,-0.0234375,-0.046875,-0.0234375,0.03125,-0.0390625,-0.078125,-0.015625,0,-0.0078125,-0.03125,-0.0078125,-0.03125,0.0625,0.015625,-0.015625,-0.109375,0.0234375,-0.015625,0.0234375,0,-0.0078125,-0.09375,-0.015625,-0.0546875,-0.0625,0.015625,0.03125,-0.0625,0.0625,-0.0859375,0.0390625,-0.046875,-0.0078125,-0.015625,-0.0078125,-0.015625,-0.0234375,0.03125,0.125,-0.0703125,-0.0078125,-0.0625,-0.015625,-0.0234375,0,-0.046875,-0.0234375,-0.015625,0.0390625,-0.0234375,0.0234375,0.015625,0.015625,-0.0234375,-0.015625,0.0078125,-0.0078125,0.0078125,0,0,0.0078125,0,0.015625,0.015625,-0.015625,-0.0625,0.03125,-0.078125,-0.0390625,0.0703125,0.0078125,-0.03125,-0.0234375,0.03125,-0.03125,0.0234375,0.0078125,-0.046875,0.0703125,-0.015625,-0.0078125,0.0078125,0,0.0234375,0,-0.046875,0.03125,0.078125,-0.0234375,0,-0.046875,0,0,-0.015625,0.0078125,0,0.0078125,-0.0078125,-0.0078125,-0.0078125,0.0625,-0.0546875,0.09375,-0.0625,-0.0859375,0.0234375,-0.03125,-0.046875,-0.0078125,0.0078125,0.0390625,0.0546875,-0.015625,0.0078125,0.03125,-0.0078125,-0.0234375,0.0078125,-0.0078125,0.0859375,0.015625,-0.0390625,0.0234375,-0.109375,-0.03125,-0.046875,-0.0234375,0.03125,-0.03125,0,-0.0078125,0.0234375,-0.0078125,-0.015625,-0.0390625,0,0.0625,-0.03125,-0.0703125,-0.0078125,0.0078125,0.015625,0.0078125,-0.0234375,0.0078125,-0.0234375,0.015625,0.03125,-0.046875,-0.0234375,-0.0234375,0.0078125,0,0,0.015625,0,-0.015625,0.0078125,-0.015625,-0.0234375,0,0,-0.0078125,-0.015625,0.046875,-0.0625,-0.0078125,-0.015625,-0.046875,0,0.0234375,0.0234375,0.03125,-0.0078125,-0.0625,0.0078125,0.0234375,0.03125,0,-0.03125,-0.015625,-0.03125,0.0859375,-0.015625,-0.078125,0.03125,-0.03125,-0.0234375,-0.0234375,-0.015625,-0.015625,0.015625,-0.015625,0,0.0078125,0.0234375,-0.0078125,0,0,0,-0.0078125,0.0078125,-0.0625,-0.0390625,0.0546875,0.015625,-0.0234375,0.0234375,0.0390625,-0.0703125,0,0.03125,-0.03125,0.0078125,-0.0078125,-0.015625,0,0.0078125,0.0390625,0.0625,-0.0234375,0.0390625,-0.0546875,-0.0234375,0.0078125,-0.0078125,-0.015625,0.03125,0,-0.0078125,-0.046875,0,-0.0078125,0.0078125,0.03125,-0.0703125,-0.046875,0,-0.0703125,0.0390625,0.046875,0.0234375,0.015625,-0.015625,0.015625,0.0703125,0.046875,0.0234375,-0.046875,-0.0078125,-0.0234375,-0.0078125,-0.0078125,-0.0390625,0.0078125,-0.0625,0.0234375,-0.03125,-0.0234375,0.015625,-0.015625,0.0078125,-0.0546875,0.0234375,-0.0234375,-0.0234375,-0.0078125,0.0390625,-0.015625,0,0.03125,-0.03125,0.046875,-0.0546875,-0.0078125,0,-0.0546875,0.0234375,0.0078125,0,0,-0.015625,-0.015625,-0.0078125,0.078125,-0.0234375,0.0078125,-0.0078125,-0.0390625,0.078125,0.0546875,0.0078125,0.015625,-0.0859375,-0.078125,-0.0078125,-0.0390625,0,0.0078125,-0.078125,-0.03125,0.03125,0.09375,0.03125,-0.0234375,0.0234375,0,0.015625,-0.0859375,-0.0390625,-0.0390625,-0.0390625,0.03125,0.0078125,-0.0078125,-0.0234375,0,0.0234375,0.0234375,-0.03125,-0.0078125,0.0625,0.015625,-0.0234375,0,0.0859375,-0.0234375,0.0390625,0.0078125,-0.015625,0.0078125,0.0078125,-0.015625,0,-0.0390625,-0.0546875,-0.03125,-0.0078125,-0.046875,0.09375,-0.0234375,-0.0078125,0.0078125,-0.0078125,0,-0.0078125,0,0.0078125,0.0078125,0.015625,-0.0078125,0.0234375,-0.0625,0.03125,0.03125,-0.0078125,0.046875,-0.015625,-0.015625,0,0,-0.046875,-0.03125,0.0078125,0.0078125,0.078125,0.046875,-0.0078125,0,0,-0.0078125,-0.015625,-0.0390625,0,-0.0234375,-0.0234375,0.015625,0.0625,-0.0234375,0,0.0078125,-0.015625,0.015625,-0.015625,0,0,-0.0078125,-0.0078125,-0.0390625,0.03125,-0.03125,-0.0234375,-0.0703125,-0.0390625,-0.0234375,-0.0078125,0.03125,-0.0390625,0.015625,-0.0625,-0.015625,-0.0390625,0.0859375,-0.03125,-0.0703125,-0.046875,-0.0078125,-0.0625,-0.0078125,-0.015625,0,-0.0390625,-0.0625,-0.015625,-0.0859375,0,0.015625,-0.0078125,-0.0390625,-0.0546875,-0.0703125,-0.0234375,0.0078125,-0.0390625,-0.0234375,-0.0859375,-0.0546875,-0.046875,-0.015625,-0.03125,0.0078125,0.015625,0.0390625,0.0078125,-0.0078125,-0.015625,0.046875,0,-0.03125,0.0078125,-0.0546875,0.03125,0.0234375,0.078125,0.0078125,0,-0.0234375,-0.0234375,-0.0078125,0.0078125,0.0078125,0,0.0234375,-0.0234375,0.015625,-0.0390625,-0.0390625,-0.0234375,0.015625,-0.0078125,-0.03125,-0.046875,-0.03125,-0.0234375,-0.078125,0.078125,-0.0078125,-0.0078125,-0.03125,-0.0078125,-0.0234375,-0.0859375,-0.0546875,-0.0234375,0.0234375,0,0.03125,-0.0234375,0.0078125,0,0.015625,0.015625,0,0,-0.015625,0,0.015625,-0.0078125,0.0546875,-0.03125,0.015625,0.0390625,-0.0078125,-0.0234375,0.0078125,0.0078125,0,0.03125,0,-0.015625,-0.015625,-0.0390625,0,0.0546875,0.0078125,-0.0078125,-0.03125,0.03125,0.0390625,0.0390625,0.015625,0.015625,-0.03125,-0.0234375,0.0546875,-0.0546875,0.0390625,-0.046875,-0.0625,0.0234375,-0.0234375,-0.0546875,0.015625,-0.0078125,0.1015625,-0.0078125,0.0078125,-0.0078125,-0.046875,0.0234375,0.0625,-0.0859375,0,0.09375,0.0390625,-0.03125,0.0234375,-0.0625,-0.0234375,0.0078125,-0.0234375,0,0.09375,-0.0234375,0,-0.0078125,0.0078125,0,0.0234375,0.0234375,0,-0.0234375,0.0078125,0,-0.0078125,-0.0078125,0.0234375,-0.0078125,0.03125,0.0390625,0.03125,-0.0390625,0.0390625,-0.0078125,-0.015625,-0.0078125,-0.015625,0.0234375,-0.0234375,0.1015625,-0.0234375,-0.0078125,0.046875,0.03125,0.0390625,0,0.0234375,-0.03125,0.0546875,-0.0390625,-0.078125,-0.0625,0.015625,-0.03125,0.0078125,0.03125,-0.0234375,-0.0078125,0.0390625,-0.0234375,-0.046875,0.015625,0.0234375,-0.0078125,0.0546875,-0.0390625,0.15625,-0.0390625,-0.015625,-0.0234375,-0.0546875,-0.0234375,0.1015625,0.0546875,-0.03125,0.015625,-0.0234375,-0.0078125,-0.03125,-0.015625,-0.0078125,-0.015625,0.0234375,-0.0234375,0.015625,-0.0546875,-0.03125,0.015625,0.046875,-0.0390625,0,-0.015625,-0.03125,-0.046875,-0.03125,-0.0078125,-0.015625,0.015625,0.0625,0.0546875,-0.03125,0.0078125,-0.0078125,-0.015625,-0.0078125,-0.0078125,-0.0078125,0,0,-0.0078125,-0.046875,0.0234375,0.046875,-0.0625,-0.0546875,0.0078125,0.03125,0.09375,-0.09375,0.015625,-0.0546875,0.0546875,0.015625,-0.0078125,-0.0234375,0.0625,0.0859375,-0.0390625,0.1015625,0.0078125,0.0390625,-0.0703125,-0.0078125,-0.0390625,-0.046875,0.0078125,-0.0234375,-0.0078125,-0.0078125,0.015625,0,-0.0078125,0,-0.0078125,0,-0.0078125,0.0625,-0.046875,-0.0078125,0.140625,0,-0.0625,0.078125,0.0078125,0.015625,0.0703125,0.03125,0.0703125,0.0078125,0.0078125,-0.0390625,0,-0.015625,-0.0078125,0.0078125,-0.0625,0,-0.0234375,-0.03125,-0.0625,0.046875,0.0078125,-0.03125,0,0.015625,-0.015625,0.0625,0.046875,0.0078125,-0.0390625,-0.03125,-0.0078125,0.0234375,-0.0234375,-0.015625,-0.0078125,-0.03125,0.0078125,-0.015625,-0.078125,-0.015625,0.0234375,-0.0234375,-0.03125,-0.0625,0,0.0390625,0.0234375,-0.015625,0.0078125,0.03125,0.0546875,0.03125,-0.0234375,0.015625,0.015625,-0.015625,-0.015625,0.015625,0,-0.015625,0.0234375,-0.0546875,-0.015625,0.0078125,-0.0234375,0.015625,-0.015625,0.046875,0.015625,-0.015625,0.0234375,-0.0546875,-0.03125,-0.0078125,-0.0546875,-0.0546875,0.0703125,0.125,-0.078125,-0.015625,-0.09375,-0.015625,-0.0625,0,-0.078125,-0.0078125,-0.015625,0.0078125,0.0078125,-0.015625,-0.0078125,-0.015625,0,0,0.015625,0,-0.015625,-0.0078125,-0.0546875,0.015625,0.0625,-0.0234375,-0.03125,-0.0078125,-0.0234375,-0.0078125,-0.0078125,0.0234375,0.0390625,0,0.0390625,-0.03125,-0.0078125,0.0390625,0.0390625,0.046875,-0.03125,-0.0390625,-0.0234375,0.015625,-0.0234375,0,-0.015625,0.0234375,0,-0.0234375,0.015625,-0.03125,-0.03125,0.015625,-0.03125,0.0625,0.0078125,0.03125,-0.0546875,-0.0234375,-0.015625,-0.0546875,0.0390625,0,-0.0078125,0.0390625,-0.0390625,-0.046875,0,0.0625,0.09375,0,0.0546875,-0.0390625,0.03125,-0.0546875,-0.0625,0.078125,0,0.0078125,-0.0078125,0,-0.0078125,-0.046875,0,-0.046875,0,0.0390625,-0.0390625,-0.0234375,-0.0390625,-0.0546875,0,-0.0390625,0.0625,0.015625,-0.03125,0,0.0703125,-0.0078125,0.0859375,0.03125,-0.0234375,-0.0234375,-0.0703125,0.046875,0.0546875,0.03125,0.0234375,-0.0078125,-0.0625,0.0078125,-0.09375,0.015625,0.0078125,-0.0234375,0.0078125,0.1484375,-0.015625,-0.0078125,-0.0234375,-0.0703125,-0.046875,-0.0390625,-0.046875,-0.078125,-0.03125,0,0,-0.0078125,-0.03125,-0.015625,-0.046875,0,0,0.046875,0.1328125,0.0546875,-0.109375,0.0234375,-0.015625,0,-0.015625,-0.03125,-0.015625,-0.0546875,-0.0234375,-0.046875,-0.0234375,-0.0234375,0,-0.015625,0,0.0078125,0.0234375,0.0078125,0.0078125,-0.0703125,0,-0.015625,0.0078125,0.0859375,0,0,-0.0078125,-0.015625,0.0078125,0.0078125,-0.0078125,0,0,0.015625,-0.0234375,-0.015625,-0.0078125,0.0234375,0.046875,0,-0.0078125,-0.0234375,-0.0078125,0.0234375,0,0,0.0078125,0,-0.0078125,-0.0234375,-0.0234375,-0.0234375,-0.0625,-0.0078125,-0.0390625,0.046875,0.0546875,-0.0234375,-0.0390625,-0.046875,0.0078125,-0.0078125,-0.0078125,0,-0.0078125,-0.0078125,-0.0078125,0.0078125,0.0078125,-0.03125,0.0234375,0.03125,-0.0390625,-0.03125,-0.078125,0,-0.0390625,0.015625,-0.015625,0.078125,-0.046875,-0.0234375,0.0234375,0.015625,-0.0234375,0.046875,-0.015625,0.015625,0.078125,0,-0.0546875,-0.0078125,0.0546875,-0.0390625,-0.046875,-0.078125,0.0390625,0.03125,0.0078125,0.03125,-0.03125,0,-0.015625,-0.03125,-0.0234375,-0.015625,0.0078125,0.046875,-0.03125,0,-0.015625,-0.0234375,-0.0234375,-0.0234375,-0.03125,-0.0234375,-0.0234375,-0.015625,0.03125,-0.0078125,-0.0078125,-0.015625,-0.015625,-0.0234375,-0.015625,-0.015625,-0.015625,-0.03125,0.0078125,0.0078125,0.0078125,-0.0078125,-0.0234375,0,0.015625,0,0.015625,0.03125,-0.015625,0.015625,-0.0234375,0,-0.03125,0.0390625,-0.0078125,-0.0078125,-0.0390625,-0.0078125,-0.0234375,-0.0078125,-0.015625,-0.015625,-0.0078125,-0.015625,-0.0078125,-0.0078125,-0.03125,0,0.0390625,-0.0078125,0.015625,0,-0.0078125,0,0.0078125,-0.0078125,0.0234375,0.0078125,-0.03125,-0.046875,0.0078125,-0.0078125,0.015625,0.015625,0,-0.0078125,0.015625,0.015625,0,-0.0234375,-0.0078125,0.0234375,0.0078125,-0.015625,-0.015625,-0.0234375,0.03125,0.0703125,0.0234375,-0.03125,0.0078125,0.0859375,-0.015625,-0.0390625,-0.078125,-0.0546875,-0.015625,-0.0546875,0,0.0546875,0.0390625,-0.015625,-0.0234375,0.0546875,-0.015625,0.0078125,0.0078125,-0.0078125,-0.0859375,0.0546875,0.0078125,-0.03125,-0.0390625,0.015625,0,-0.03125,-0.0234375,0.0390625,0.015625,-0.0234375,-0.0234375,-0.015625,0.015625,-0.0234375,-0.015625,0.0078125,-0.0078125,0.0546875,-0.015625,0.0390625,-0.0625,-0.0234375,0.0078125,0,-0.015625,0.046875,0.0546875,-0.0078125,-0.0546875,-0.015625,-0.046875,0.015625,-0.046875,-0.0234375,0.0703125,-0.03125,-0.0078125,-0.03125,-0.015625,0,-0.0078125,-0.015625,-0.078125,-0.09375,-0.0546875,-0.0078125,-0.0078125,0.046875,0.0078125,-0.0703125,-0.0703125,-0.015625,0.0390625,0.0390625,-0.0078125,-0.0625,-0.046875,-0.0078125,-0.0078125,-0.0390625,0,0.046875,-0.046875,-0.0078125,-0.015625,-0.0078125,-0.0546875,-0.03125,-0.015625,-0.0234375,-0.03125,-0.09375,-0.0078125,-0.0390625,0.0390625,-0.0078125,-0.0703125,-0.0703125,-0.0390625,0.03125,-0.0078125,-0.0234375,0.015625,0.15625,-0.0234375,0,-0.03125,-0.0234375,0.015625,-0.0234375,-0.0234375,0.0390625,-0.0390625,0.0234375,-0.03125,-0.0390625,0.0078125,0,-0.015625,0.0390625,0.09375,-0.0078125,0.0078125,-0.015625,0,0,0,-0.0234375,0,-0.0078125,0,-0.015625,0.0625,-0.046875,-0.0546875,-0.1015625,-0.078125,-0.0078125,0.1015625,0.0234375,0.0078125,0.078125,-0.0234375,0.03125,-0.03125,-0.015625,0.0390625,-0.015625,-0.03125,0.03125,-0.0078125,0.03125,-0.0703125,-0.0234375,-0.046875,-0.078125,0.0078125,0.03125,0,-0.015625,-0.0078125,-0.0078125,0,0.0078125,0.0078125,0,0.0078125,0.0234375,0.0078125,0.0390625,0.03125,0.03125,-0.03125,-0.0625,0.0546875,0,0.0078125,0.1484375,-0.0625,-0.0078125,-0.09375,-0.078125,0.015625,0.0078125,-0.03125,0.015625,-0.0078125,0.0078125,0.0078125,-0.0078125,0.015625,0.015625,-0.0078125,0.0078125,0.0234375,0,0.0078125,0.015625,0.0078125,0.0546875,0.0234375,-0.03125,0.0234375,0,-0.0234375,0.0546875,0,0.015625,-0.015625,-0.0625,0.015625,-0.0390625,-0.015625,0.015625,0.0234375,0,0.0078125,-0.0078125,-0.0234375,-0.03125,-0.0625,0,0.0703125,0.0078125,-0.0390625,-0.0234375,-0.0390625,-0.03125,-0.0078125,-0.015625,0.0078125,-0.015625,-0.015625,0.03125,-0.03125,-0.0078125,-0.046875,-0.0390625,-0.015625,-0.015625,-0.0234375,0,0.0078125,0.109375,0.0390625,-0.0078125,-0.0390625,0,0.0546875,0.046875,0.0078125,-0.0078125,-0.0234375,-0.015625,0.0078125,0,0.0078125,0.0078125,0,0.0078125,0,-0.0234375,-0.0078125,0.0078125,0.0078125,0.015625,0,0.125,-0.015625,-0.03125,0.046875,-0.0390625,-0.0078125,0.03125,0,-0.0390625,0.0625,-0.015625,-0.0234375,-0.0234375,0,-0.03125,-0.0390625,-0.0078125,-0.046875,-0.125,0.0234375,-0.0234375,0.03125,-0.03125,0.0390625,0.0703125,0.0546875,0.0234375,-0.03125,0.0703125,-0.03125,-0.0859375,-0.0859375,-0.0390625,-0.09375,-0.015625,-0.046875,-0.015625,-0.078125,-0.046875,-0.046875,-0.0546875,-0.0078125,0,-0.0234375,0,-0.0078125,-0.0234375,-0.0703125,-0.0234375,0.0390625,-0.015625,-0.03125,0.015625,-0.0078125,0.03125,-0.046875,-0.03125,-0.0859375,0,0.03125,-0.046875,-0.03125,0.0390625,-0.0390625,0.03125,-0.0390625,0.03125,-0.03125,0,-0.0078125,-0.0703125,-0.0078125,-0.0703125,-0.015625,-0.0546875,-0.0078125,-0.078125,0.0078125,-0.0703125,-0.0859375,0.046875,-0.015625,0.0078125,-0.0234375,-0.046875,-0.0234375,0.0234375,0.015625,0.0078125,-0.046875,0.1015625,-0.03125,0.0078125,-0.0234375,-0.0078125,-0.015625,-0.078125,-0.0234375,0.0078125,-0.078125,0.015625,0.0546875,0.0546875,0,-0.078125,-0.078125,-0.0625,-0.046875,0.0546875,-0.03125,-0.015625,-0.03125,0.0078125,-0.0546875,-0.109375,0.0078125,0.0546875,0.0234375,0.046875,-0.03125,-0.0859375,-0.03125,-0.0234375,-0.015625,-0.0390625,-0.03125,0.0859375,-0.0390625,-0.0234375,-0.0859375,0,-0.015625,0.0234375,0,-0.015625,-0.078125,0.046875,0.0078125,-0.015625,0.0625,0.046875,0.015625,-0.0234375,0.015625,0.0078125,0,0,-0.0078125,0.015625,-0.0078125,-0.0234375,-0.0234375,-0.015625,-0.03125,-0.0546875,-0.0078125,0.03125,-0.1015625,0.0625,0.0234375,-0.0234375,-0.0078125,-0.03125,-0.0390625,0.1015625,-0.0546875,-0.0546875,0.0234375,-0.0234375,-0.0546875,0.0078125,0,-0.015625,-0.0859375,-0.0625,0.0859375,-0.0390625,-0.0625,-0.046875,0,-0.015625,0.0078125,-0.0078125,0.0078125,-0.015625,-0.015625,-0.0078125,0,0,0.0234375,0.015625,-0.015625,0,-0.046875,-0.03125,0.0078125,-0.046875,0.015625,-0.0546875,0.078125,-0.015625,-0.046875,0.09375,-0.0234375,-0.0859375,0.03125,-0.0078125,-0.0859375,0.015625,-0.03125,-0.015625,0.03125,-0.046875,0.0078125,-0.03125,0.015625,-0.0078125,0.046875,-0.015625,0.015625,-0.03125,0.03125,0.03125,0.0390625,0.078125,0.0703125,0.078125,-0.0234375,-0.03125,0,0,0.015625,0,-0.0078125,0,0,0.0078125,0.0234375,0.09375,-0.0234375,-0.015625,0.0078125,-0.015625,-0.0234375,0.0078125,0.0078125,0.046875,0.0078125,-0.015625,0.0078125,0.0078125,0.0234375,0.015625,-0.015625,0.0078125,0.0078125,-0.0234375,-0.0234375,0,0.03125,-0.0234375,-0.03125,0.125,0.078125,-0.046875,-0.03125,0.03125,-0.0078125,0.015625,0.0078125,0.0234375,0.0078125,-0.015625,-0.0078125,0.046875,-0.0078125,-0.0234375,-0.03125,-0.015625,-0.015625,-0.0078125,0.0078125,-0.03125,0.0078125,0.0078125,-0.0078125,0,0.0078125,-0.0546875,0.03125,-0.0078125,0.03125,0.0625,0,0.0625,-0.046875,0.078125,-0.0234375,-0.015625,-0.0234375,0.015625,-0.03125,0.0390625,0.0234375,0.03125,0.03125,0.015625,0.0234375,-0.0390625,-0.078125,0.0234375,-0.015625,-0.0078125,0.09375,0.0078125,-0.0390625,-0.03125,-0.125,0.0546875,-0.046875,0.046875,0.0546875,0.0234375,0,0,-0.046875,-0.0625,-0.0234375,0.078125,0,-0.0234375,0.015625,-0.0703125,-0.078125,-0.03125,0.0390625,0.015625,0,0.046875,-0.0703125,0.0703125,0.0703125,0.140625,-0.0703125,-0.0703125,-0.0703125,-0.140625,0.0703125,-0.0234375,0.0390625,-0.0234375,-0.0546875,0.0234375,-0.0390625,0,0.1015625,0.0390625,-0.03125,-0.03125,-0.078125,-0.0234375,-0.0078125,-0.0234375,0.125,-0.0703125,0.03125,-0.09375,-0.078125,0.0625,0.0390625,-0.0703125,-0.046875,0.0078125,0.0078125,0.015625,0.0234375,-0.046875,0.0625,0.0390625,0.1171875,-0.046875,-0.0546875,-0.0625,-0.015625,0.078125,0.0546875,0.1015625,-0.0078125,0.046875,-0.0390625,-0.0078125,0.0078125,0.0703125,0.0078125,0.078125,0.046875,0.0625,-0.0234375,0.015625,-0.0234375,0,-0.0625,-0.0390625,-0.015625,-0.03125,-0.0078125,-0.0546875,0,0.0703125,-0.0390625,-0.015625,-0.046875,-0.0390625,0.0390625,0.0078125,0.015625,-0.03125,-0.0234375,-0.0390625,0.0546875,-0.0546875,-0.0234375,0.0078125,-0.046875,-0.0234375,0,-0.046875,-0.0234375,0.078125,0.0234375,0.0234375,0.015625,-0.0078125,-0.015625,0,0.0078125,-0.0078125,0,-0.0078125,0,-0.0078125,0.15625,-0.0234375,-0.046875,-0.0625,-0.03125,0,-0.0078125,0.015625,0.0390625,-0.0078125,0.0078125,0,-0.046875,-0.046875,0,-0.015625,0.03125,0.015625,0,-0.03125,0,-0.0546875,-0.1015625,-0.0546875,0.0703125,-0.0390625,0.0078125,0,0,0,0.0078125,0,0.0078125,0.015625,0.0078125,-0.0234375,0.03125,0.0234375,-0.046875,-0.03125,-0.078125,-0.0546875,0.03125,-0.0078125,0,0.046875,0.0234375,0.03125,-0.0546875,-0.0546875,0.046875,0.0078125,0.0234375,-0.0390625,0,-0.0390625,-0.0546875,0.0859375,0.109375,0.078125,-0.03125,0.0546875,-0.015625,0.015625,0.03125,-0.0078125,0,0.015625,0.03125,-0.046875,-0.0234375,0.0390625,-0.015625,0.078125,-0.0859375,-0.0703125,0.046875,0.046875,0.0234375,-0.015625,0.0078125,-0.0859375,-0.0546875,0,0.03125,0.015625,0.0078125,0.0546875,0.0546875,-0.015625,0.0390625,-0.0390625,-0.0078125,0.0078125,0.015625,-0.0078125,0,0.015625,-0.0390625,0,-0.0390625,0.015625,0.0078125,-0.0234375,-0.0234375,0,-0.015625,0.046875,-0.0234375,0.03125,0.0078125,0.0703125,-0.0078125,-0.0078125,0,0.03125,0.0625,-0.046875,0.078125,0.0078125,0.0078125,-0.015625,-0.0234375,-0.09375,-0.046875,0,0,0,0.0078125,0,0.0078125,-0.015625,0,-0.015625,0.0078125,0.03125,-0.078125,-0.0390625,-0.0234375,0,0,0,-0.0078125,0.0390625,0.03125,-0.03125,0,0.03125,-0.078125,0.015625,-0.0390625,-0.0703125,-0.046875,-0.109375,-0.015625,0.0859375,-0.046875,0,-0.015625,0,0.0859375,-0.0234375,0.0390625,0.140625,-0.046875,0.0078125,-0.0703125,-0.0703125,-0.0703125,-0.09375,0.1328125,0.0625,-0.078125,0.0078125,-0.140625,-0.03125,0.1015625,-0.046875,-0.140625,0.046875,0,-0.0234375,-0.015625,-0.0234375,-0.0390625,-0.0859375,0,0.015625,-0.046875,0.0234375,0.0234375,-0.0234375,-0.0234375,0,0.015625,0.03125,-0.0078125,0.0625,-0.03125,0.0078125,0,-0.0625,0.046875,0.0078125,0.0390625,0.0546875,-0.0078125,-0.015625,0.015625,0.03125,0,-0.0078125,0.046875,-0.03125,0.0859375,-0.0546875,-0.03125,-0.0234375,-0.078125,-0.078125,-0.0234375,0.0078125,0.0703125,0.03125,-0.1015625,0,0.0078125,0.0078125,0,-0.015625,-0.015625,-0.0546875,0.046875,-0.015625,0.0703125,0.0703125,-0.03125,-0.0390625,-0.0546875,0.0546875,-0.0234375,0.015625,0.0546875,0.0234375,-0.0078125,0.09375,-0.0625,0.0078125,0.03125,-0.046875,0.109375,0.0390625,0.015625,0.0546875,-0.03125,-0.078125,-0.015625,-0.0546875,-0.0078125,0.0234375,0.0703125,-0.0078125,-0.0546875,0.03125,-0.015625,0.0078125,0,0.0859375,0.078125,0.0078125,0.015625,0,0.0078125,0.046875,0.015625,0.0234375,0.0234375,0.03125,-0.0078125,-0.0078125,0,-0.015625,-0.0078125,0.0078125,0,0.015625,0.015625,-0.015625,0.0234375,0.0234375,-0.0078125,0.0546875,0,0.0078125,-0.03125,-0.0234375,-0.0234375,-0.015625,0.0078125,0.0078125,0.015625,0.03125,0.0078125,0.0078125,0,-0.015625,-0.015625,-0.0625,0.015625,-0.046875,-0.0390625,0,0.0390625,-0.015625,-0.015625,0,-0.015625,0,0.015625,-0.0078125,-0.0078125,0,-0.0078125,0.015625,-0.0390625,-0.015625,0.015625,-0.015625,0,0.015625,-0.046875,0.078125,-0.0546875,-0.03125,-0.0078125,0.03125,0.0390625,-0.0078125,-0.0078125,0.0703125,-0.0546875,-0.03125,-0.015625,-0.0234375,0.015625,0.015625,-0.0078125,-0.046875,-0.0390625,0.015625,-0.015625,-0.015625,-0.015625,0.0390625,0.046875,-0.0234375,0,0,-0.0234375,0.03125,-0.015625,0.015625,-0.015625,0.0234375,0.0078125,-0.0078125,0.0546875,-0.015625,0,-0.015625,0.015625,-0.0234375,-0.03125,0.03125,0.015625,-0.0234375,0.03125,0,-0.0078125,-0.0078125,0.015625,0.0078125,-0.015625,0.0078125,0,-0.015625,-0.0078125,0,0.0234375,-0.015625,-0.0390625,-0.015625,-0.0390625,-0.03125,-0.0078125,-0.015625,-0.0234375,-0.03125,-0.03125,0.0078125,0,-0.03125,0.0625,0.0234375,-0.0078125,-0.03125,-0.0390625,0,-0.015625,-0.015625,-0.03125,0,0.0078125,0.0078125,-0.0078125,0.0078125,0.0078125,-0.0078125,-0.015625,0.0078125,0.0078125,-0.015625,-0.0078125,0.015625,0.0390625,0.015625,0.0078125,0,0.0703125,0.0078125,0.0078125,0,-0.0234375,-0.03125,0.0390625,-0.078125,-0.03125,-0.0234375,-0.03125,-0.03125,-0.0078125,-0.015625,-0.03125,0.0234375,-0.0625,-0.0546875,0.03125,0.0234375,0.015625,0.03125,-0.03125,-0.046875,-0.015625,-0.1015625,-0.0078125,-0.0234375,0.046875,0,0,0.015625,0.015625,-0.015625,-0.015625,-0.0546875,0.0546875,-0.0234375,0.0078125,0.0234375,0.015625,0.0078125,0.015625,-0.0234375,0.078125,-0.015625,-0.0234375,0.0234375,-0.015625,0.0234375,0,0.046875,-0.0546875,0.015625,0.0234375,-0.078125,-0.03125,0,0.0078125,0.0078125,-0.03125,0.0078125,-0.015625,0.0234375,-0.0234375,-0.015625,0.0078125,0.0078125,0.0625,0.015625,0.0625,0.0859375,-0.03125,-0.015625,-0.03125,-0.046875,-0.0078125,-0.0078125,-0.015625,-0.0546875,-0.03125,0.0234375,-0.0390625,-0.046875,-0.0625,0.0390625,0,-0.046875,-0.015625,-0.125,-0.0390625,0.015625,0,0.0078125,-0.0390625,-0.03125,0.0078125,-0.1015625,-0.015625,0.0078125,-0.015625,0,-0.0234375,0.015625,0.015625,0.0703125,0,0,-0.015625,-0.03125,-0.03125,0.0546875,-0.0234375,-0.0234375,0.1015625,-0.0078125,0.09375,0.0078125,0,-0.015625,0,-0.0078125,0.0078125,0.0390625,0.0078125,0,-0.046875,-0.03125,-0.0078125,0.0390625,0.0546875,0.0078125,-0.0234375,0,-0.015625,-0.015625,-0.0390625,-0.015625,0.0078125,-0.0078125,-0.0078125,0.0234375,-0.015625,0.0078125,0,0,0.015625,-0.0234375,0.09375,0.109375,-0.0703125,-0.0859375,0.03125,-0.0234375,-0.0078125,-0.0234375,-0.0546875,-0.1328125,-0.0390625,0.0390625,-0.0390625,0.0703125,-0.03125,0.0859375,-0.046875,-0.03125,0.0234375,-0.0546875,0.0625,0.0546875,-0.046875,0.0234375,-0.015625,-0.0625,0.0234375,-0.0078125,0.0078125,-0.0078125,0,0,0,0,0,0.03125,0.0625,-0.09375,0.0078125,-0.109375,-0.0078125,-0.0546875,0.015625,-0.0625,0.0234375,-0.0234375,0.0390625,-0.1015625,-0.0546875,0.015625,0.03125,-0.0078125,0.046875,-0.0703125,-0.015625,0.109375,-0.09375,-0.015625,0.109375,-0.09375,-0.015625,-0.0234375,0.015625,0.03125,0.1015625,-0.046875,0.0078125,0.0234375,-0.0078125,0.015625,-0.0078125,-0.0390625,-0.0546875,-0.015625,-0.0078125,0.015625,-0.0703125,-0.0390625,0.03125,-0.015625,0,-0.046875,0,0.046875,-0.03125,-0.0234375,-0.015625,-0.0234375,0.0859375,0.015625,0.03125,-0.015625,-0.0703125,-0.0390625,0.0703125,0.03125,-0.015625,-0.03125,-0.046875,0.0390625,-0.0078125,-0.03125,-0.0390625,0.03125,0.0234375,0.046875,-0.0234375,-0.0390625,-0.015625,0.015625,0,-0.015625,-0.0390625,-0.0703125,0.015625,0,-0.03125,-0.03125,0.0546875,-0.046875,-0.046875,0.0390625,0.015625,0.03125,0,-0.015625,-0.0078125,-0.015625,-0.0078125,0.0078125,0.0078125,0.015625,-0.015625,0.0078125,-0.0546875,0.0625,-0.015625,0.0390625,-0.0078125,0.0234375,-0.03125,0.015625,-0.03125,-0.046875,0,0,0.0390625,0.015625,0.046875,-0.0390625,-0.0625,0.015625,0.046875,0.0390625,0.0234375,0.0390625,0.0078125,-0.125,0.078125,0.03125,0.0390625,0.09375,0.0234375,-0.078125,0.0546875,-0.015625,-0.03125,0.0234375,0.015625,0.0234375,0.078125,0,-0.0234375,0.015625,0.0390625,-0.0625,0.109375,0.0234375,0.03125,0.09375,0.0078125,-0.078125,0.0078125,-0.0390625,-0.0625,-0.03125,-0.0390625,0.046875,-0.0546875,0.0234375,-0.1328125,0.0078125,0.140625,-0.015625,-0.0859375,-0.0234375,0.140625,0.03125,0.03125,-0.03125,0.0390625,-0.015625,-0.0703125,0.0234375,-0.078125,0.0546875,-0.03125,-0.0390625,0.0234375,-0.0546875,0.03125,0.03125,-0.0234375,0,-0.015625,-0.0390625,0.0078125,0.0390625,-0.09375,-0.0625,0.0390625,0.015625,-0.0078125,-0.0390625,-0.0546875,0.0625,0.015625,-0.140625,0.0546875,0.046875,0.0234375,0.109375,-0.0703125,-0.0234375,0.078125,-0.0078125,0.015625,0.0859375,-0.0234375,-0.015625,-0.046875,-0.125,0.046875,-0.03125,-0.0625,-0.0546875,0.03125,-0.03125,0.0234375,-0.0078125,-0.03125,0.078125,0.0390625,-0.0546875,0.0703125,-0.078125,-0.015625,-0.03125,0.0078125,0.0546875,0.0234375,0.078125,-0.0546875,-0.0078125,0.0234375,-0.0625,0,-0.09375,0.0859375,-0.0234375,-0.046875,-0.015625,-0.0625,-0.0625,-0.03125,-0.015625,-0.0390625,0,-0.015625,-0.0078125,0,0.0078125,0.0078125,0,0.015625,0.0078125,-0.0078125,0.0703125,0.125,0.0234375,-0.0078125,-0.0546875,0.0078125,0,-0.0703125,0.03125,-0.046875,0.046875,-0.0703125,0,-0.078125,0,-0.015625,-0.0625,0.0703125,-0.03125,0.03125,0.0234375,0.0859375,-0.03125,0.0703125,0,0.0078125,0.0546875,-0.0078125,0,-0.015625,0,0.0078125,0.015625,0,0.0078125,-0.0078125,-0.015625,-0.046875,-0.015625,0.0078125,0.015625,-0.046875,0.125,0.1015625,-0.0234375,-0.0546875,-0.0078125,-0.0390625,0,0.015625,0,-0.0390625,-0.0546875,0.0078125,0,0.015625,0.0546875,-0.046875,-0.109375,0.015625,0.046875,-0.0078125,0.0390625,-0.0078125,0.0078125,0.0234375,0.03125,0,0.0078125,0.0390625,0.03125,0.015625,0,-0.015625,0.0625,-0.0078125,0,-0.03125,0.03125,0.0703125,-0.0390625,0.015625,-0.0546875,-0.0234375,0.0078125,-0.0234375,0.0234375,0.03125,0.015625,-0.03125,-0.0078125,-0.015625,-0.046875,0,0.0078125,0,-0.0078125,-0.0234375,0,-0.0078125,-0.0234375,-0.0078125,0,0.0078125,0.046875,0.0234375,0.0078125,0.015625,0.0078125,0.015625,0.046875,0.046875,0.1171875,-0.0234375,0.0234375,0.0234375,-0.046875,-0.0390625,0.03125,-0.03125,0.015625,0.0859375,-0.0390625,0,0.03125,-0.0390625,-0.015625,0,-0.0078125,-0.0078125,-0.0234375,0,0,-0.0234375,-0.015625,0.0390625,-0.0234375,-0.03125,-0.0078125,0.015625,0.03125,0.0078125,-0.015625,-0.0078125,-0.0390625,0.0234375,-0.0390625,-0.0625,-0.0390625,0.0234375,0.0078125,0.015625,0,0.0234375,0.0703125,0.0546875,0.015625,-0.0234375,-0.0234375,-0.03125,-0.015625,0.03125,-0.0078125,-0.0234375,-0.0546875,-0.0234375,-0.0546875,-0.0625,-0.015625,0,0.0078125,-0.015625,-0.0234375,0.015625,-0.0234375,-0.078125,0.0234375,0.03125,-0.0234375,0,0.046875,0.0078125,0.0078125,-0.0234375,-0.0390625,0.015625,-0.0546875,-0.078125,-0.0625,0,0.046875,-0.03125,0.0234375,0.046875,-0.0234375,-0.0546875,-0.09375,-0.015625,0.0625,-0.03125,0.0625,-0.0390625,-0.046875,-0.0390625,-0.0390625,0.0078125,-0.0234375,-0.0078125,0.0546875,0.0234375,-0.046875,-0.015625,-0.03125,-0.046875,-0.078125,-0.03125,-0.0390625,-0.0078125,-0.046875,0.078125,-0.0390625,0.0390625,0.03125,0.0234375,0.078125,0.09375,0.0234375,0.046875,-0.0546875,0.03125,-0.078125,0.03125,0.046875,-0.078125,0.03125,-0.0390625,-0.03125,0.0703125,-0.03125,0.046875,-0.015625,-0.03125,-0.0703125,-0.0234375,0,-0.0546875,0.015625,-0.015625,0.0078125,0.0390625,-0.078125,0.015625,-0.0625,0.0546875,-0.046875,0.0234375,0.0390625,-0.0078125,-0.0234375,-0.0234375,-0.03125,-0.0625,-0.078125,-0.0390625,-0.0078125,-0.0234375,-0.046875,-0.03125,-0.0234375,-0.0234375,-0.0234375,-0.0546875,-0.0390625,-0.015625,0,0.03125,-0.0078125,0.09375,-0.0234375,-0.015625,0,0.0234375,0.015625,0.0078125,-0.015625,0,0.015625,-0.0078125,0.0234375,0.0078125,0,-0.015625,0.078125,0.0546875,0.03125,-0.0078125,0.0234375,0.015625,0.0078125,0,0.0234375,0.03125,-0.015625,-0.0078125,-0.015625,-0.0546875,-0.0234375,0.0078125,-0.0234375,-0.0234375,-0.0390625,-0.046875,0.109375,-0.0234375,-0.03125,-0.015625,0.0078125,0,-0.015625,0,-0.0078125,0,0,-0.0078125,0,-0.0546875,-0.0078125,0.0546875,0.0234375,-0.0546875,-0.0234375,0.0546875,-0.0234375,-0.0390625,-0.0625,-0.0234375,0.0234375,-0.09375,0,0.09375,-0.046875,0.015625,0.0234375,0.0078125,0.0234375,-0.0703125,-0.1171875,0.0390625,0.1015625,-0.0546875,-0.0390625,0.0078125,0.0078125,-0.046875,-0.046875,0.0078125,0,-0.015625,-0.046875,0.015625,-0.0390625,0.0234375,0.0546875,0,0.0390625,-0.0078125,-0.0625,0.015625,-0.0078125,-0.015625,-0.015625,0.015625,0,0.0703125,-0.0234375,0.0625,-0.015625,0.0078125,-0.0234375,-0.0234375,0.0078125,-0.03125,-0.0078125,0.03125,0.03125,-0.015625,-0.015625,0.03125,-0.0078125,0,0.015625,0.015625,0.015625,0.046875,-0.0390625,-0.0078125,-0.0078125,0.015625,0,-0.046875,0.0234375,0.0546875,-0.09375,0.0078125,-0.0546875,-0.0703125,-0.0546875,-0.0078125,0,0.015625,-0.0703125,0.046875,0.015625,-0.046875,-0.0078125,0,0.0078125,-0.015625,-0.03125,-0.0078125,0,0,0.0078125,0.0078125,-0.0078125,0.0078125,0.03125,0.0078125,-0.015625,0,-0.03125,-0.0078125,0.0390625,0.09375,-0.03125,-0.0078125,0.015625,-0.0390625,-0.0390625,0.046875,0.015625,-0.015625,0,0.015625,-0.109375,-0.015625,-0.03125,0.015625,0.0859375,-0.015625,-0.0078125,0.0234375,0.03125,-0.0859375,0.171875,-0.0625,-0.0390625,-0.0078125,-0.015625,-0.046875,0.0078125,-0.046875,0.03125,0.046875,-0.0390625,-0.015625,-0.046875,-0.09375,-0.0078125,-0.0234375,-0.0234375,-0.0390625,-0.0703125,0.0078125,0.140625,0,-0.0078125,-0.046875,0.0234375,0,-0.03125,-0.0546875,-0.015625,-0.015625,-0.0546875,0.046875,-0.0234375,-0.0390625,-0.03125,-0.0625,0.046875,-0.0546875,0.0546875,-0.0546875,-0.0078125,0.0078125,0,-0.015625,-0.015625,-0.0546875,-0.0234375,0.1015625,-0.0859375,-0.0625,-0.0625,-0.0390625,-0.0078125,0.078125,-0.0390625,-0.0078125,-0.0390625,-0.0546875,-0.0078125,-0.0390625,0,-0.015625,0.0234375,0,-0.046875,0.078125,-0.0390625,0.0390625,0.0234375,0.0546875,0.0859375,-0.0546875,0.046875,-0.0859375,0.0078125,-0.078125,-0.046875,0.03125,0.0390625,0.046875,0.0625,-0.1328125,-0.015625,0.015625,-0.015625,-0.015625,-0.03125,-0.0390625,0.046875,-0.046875,-0.03125,0.015625,0.0234375,0,0,-0.015625,0.046875,0,0.0390625,-0.046875,-0.0390625,0.046875,0.0078125,-0.0078125,-0.0625,-0.0546875,-0.0234375,-0.0234375,0.0546875,0,0,0.0078125,0.015625,0.0078125,0,0.015625,-0.0078125,0,0,0.0078125,-0.015625,0,-0.046875,-0.03125,0.0546875,0.015625,-0.015625,0.015625,0,-0.0078125,-0.0390625,0,-0.0078125,0.0078125,0.015625,-0.0390625,0,-0.015625,-0.0078125,-0.015625,0.0078125,0.0234375,0.046875,0.0078125,-0.046875,0.03125,-0.0078125,-0.03125,0.03125,0.0078125,-0.0078125,0,0.0078125,-0.0078125,0,0,0,-0.0078125,-0.015625,-0.0390625,0.015625,0.015625,0.0078125,0.0078125,-0.015625,-0.0234375,-0.0234375,0.078125,0.03125,0.015625,-0.0390625,-0.0234375,-0.0234375,-0.015625,-0.015625,0.03125,0.0390625,0.046875,-0.015625,-0.0390625,-0.0078125,-0.0390625,-0.015625,0,0,0.0234375,0,-0.015625,-0.03125,0.0234375,0.015625,0,-0.0234375,-0.0078125,-0.046875,0.078125,-0.015625,0.03125,0.0078125,-0.0390625,-0.0234375,0,0.0234375,-0.0078125,0.0546875,-0.0390625,0.015625,0,0,0.0078125,-0.0234375,0,0.0078125,-0.0078125,-0.015625,0.015625,0.0078125,-0.0078125,0,-0.015625,0,0.0234375,-0.015625,0.015625,-0.015625,-0.0234375,0.0234375,0,-0.0078125,-0.0234375,0.0078125,-0.0078125,-0.046875,-0.0546875,0,-0.015625,0.0234375,0.015625,-0.0078125,-0.03125,-0.015625,-0.0546875,-0.0234375,0.0078125,0.0078125,0.015625,0.0234375,-0.0078125,-0.0078125,0.015625,0.0078125,0,-0.0078125,-0.015625,0.015625,0,0,-0.0390625,0,0.0078125,0.0234375,0.0234375,0.0234375,-0.015625,-0.015625,-0.015625,0.03125,0,0.0625,0.0234375,-0.0703125,-0.0078125,0,-0.015625,-0.0078125,0.0703125,0.1171875,-0.0546875,-0.0390625,0,-0.0546875,-0.0234375,-0.0078125,0.015625,-0.0703125,0.03125,0.0390625,-0.015625,-0.0703125,-0.015625,-0.0078125,-0.0234375,0.0078125,0.015625,0.0234375,-0.0234375,0,0.0078125,0.0078125,-0.015625,-0.0390625,0.0078125,-0.0390625,-0.0546875,-0.03125,0.0625,0,-0.0625,-0.0078125,0.015625,-0.03125,0.0625,0,0.0703125,0.0390625,-0.1015625,-0.0234375,-0.0234375,0.0234375,-0.0078125,-0.0390625,0.0546875,0,-0.03125,0.0078125,-0.078125,-0.015625,-0.0234375,-0.03125,-0.0078125,0.046875,-0.03125,0.015625,-0.0625,-0.0078125,-0.0234375,0,-0.03125,0.03125,0.0078125,0.0234375,0.0234375,0,-0.03125,-0.03125,0.0078125,0.03125,0.046875,0.03125,0.0078125,-0.0078125,0.0234375,0.03125,0,0.0078125,-0.03125,-0.078125,0.0078125,0.078125,0.0390625,-0.0546875,-0.015625,-0.015625,-0.0234375,-0.0390625,-0.0234375,0.015625,0.0546875,0.0078125,0.03125,-0.0078125,-0.0234375,-0.015625,-0.0546875,0.03125,-0.0390625,-0.046875,0.078125,-0.0546875,-0.0234375,0.0078125,0,-0.0078125,-0.046875,0.0078125,-0.015625,0.0078125,0.0234375,0.0078125,-0.015625,-0.015625,0.0234375,-0.0234375,-0.015625,-0.03125,-0.0234375,-0.03125,0,-0.015625,-0.0390625,-0.0234375,0.0078125,-0.015625,-0.0078125,0,0.0078125,-0.0078125,-0.0078125,0.0078125,0.0078125,0.0234375,-0.0234375,0,-0.0390625,-0.03125,-0.0390625,0,0.0078125,0.0078125,-0.0078125,0.0078125,0,-0.03125,0.015625,-0.0234375,0,0.0078125,-0.015625,-0.03125,0.0390625,0.015625,0.0234375,0.046875,-0.015625,-0.0234375,-0.0078125,-0.03125,0,0,-0.0078125,0.015625,0,0.015625,0,0.0078125,0.0078125,0.015625,0.0078125,0.0234375,0.046875,-0.03125,0.0078125,-0.0234375,-0.0078125,-0.015625,0.046875,0.015625,-0.0234375,-0.046875,0,-0.015625,-0.0078125,-0.0234375,0,-0.03125,0.046875,0.03125,-0.015625,0.015625,-0.015625,-0.015625,-0.0234375,-0.0390625,-0.0234375,-0.0390625,-0.0234375,0,0.0078125,-0.015625,0.0078125,0.0078125,0,0.046875,-0.0078125,0,0.0234375,-0.0703125,0.0078125,0.0234375,-0.0078125,0.0234375,0.0546875,-0.0078125,0,0.0078125,-0.015625,0.015625,0,-0.015625,0,0.015625,-0.015625,-0.0078125,0,-0.0078125,-0.0078125,0.0078125,0.0078125,0.015625,0.0234375,-0.03125,-0.0234375,-0.03125,-0.0234375,-0.0078125,0,0,0,0.0703125,-0.0234375,-0.0390625,-0.0078125,-0.03125,0,0,-0.0234375,0.0234375,-0.078125,0.015625,0.046875,-0.0078125,0.0234375,0.0078125,-0.015625,-0.0078125,0.0234375,-0.0078125,-0.0078125,0.0078125,-0.0078125,-0.0078125,-0.015625,-0.0078125,-0.015625,-0.0078125,-0.0078125,0.0078125,-0.0234375,0.0078125,-0.0078125,0,0,0,0.0078125,0.046875,0.015625,0.015625,-0.0234375,0.0078125,-0.03125,0,0.0078125,0,0.1796875,0.0234375,0.03125,-0.09375,-0.0390625,0.0078125,-0.015625,-0.0390625,-0.0234375,0.0234375,0.0546875,0.0078125,-0.046875,-0.0078125,-0.0078125,-0.0234375,0.015625,0.03125,-0.03125,-0.015625,-0.0078125,0.03125,0,0,-0.0234375,-0.0234375,0.0234375,0.015625,-0.03125,0.03125,0.0078125,0.015625,-0.015625,-0.015625,-0.0234375,-0.0078125,0.0234375,0.0234375,0.0234375,-0.0546875,-0.0078125,-0.046875,0,0.0078125,0,0.03125,0.015625,-0.015625,0.0078125,-0.046875,-0.0078125,0.015625,-0.015625,-0.0078125,0.015625,0.0390625,-0.0078125,0.0390625,0.0546875,-0.015625,0,0.0078125,-0.0078125,0.0078125,0.0078125,-0.015625,-0.015625,0,0.0078125,-0.0078125,-0.0234375,-0.0078125,0.0859375,0.0234375,-0.0234375,0.0078125,-0.0625,0,-0.0078125,0.0078125,0,0.03125,0.0234375,-0.0234375,-0.0390625,0,-0.0234375,-0.015625,0.0546875,0.0390625,-0.03125,0.03125,0,-0.046875,-0.046875,-0.0078125,0.0078125,0.0078125,0.046875,0.0078125,-0.0546875,-0.0078125,-0.03125,-0.0078125,0.0078125,-0.015625,0.015625,0.0390625,-0.03125,-0.0625,0,0,0,0.0078125,0.0234375,0,0,-0.03125,0.046875,0.0703125,-0.0625,0.0234375,0.0546875,0.03125,-0.0078125,0.0078125,-0.0078125,-0.0078125,0,-0.0078125,0.015625,0,0.0078125,0.015625,0,-0.0390625,0.0703125,0.03125,-0.0546875,0.0078125,0,0.015625,-0.046875,0.0546875,0,0.0546875,0.0078125,0.0234375,0,-0.0859375,0.0703125,-0.03125,-0.015625,0.0390625,0.015625,-0.03125,0.03125,0.015625,0.078125,-0.0234375,0.03125,0,-0.0078125,0.0078125,-0.0078125,-0.0078125,-0.015625,0,0,-0.0078125,0.0078125,0,0.046875,-0.0703125,-0.0078125,-0.015625,0,0.0234375,0.015625,-0.078125,0.0546875,-0.0078125,-0.078125,-0.0234375,0.015625,0.015625,-0.046875,-0.015625,0.015625,0.015625,0.03125,-0.0078125,0.015625,0.03125,-0.0234375,0.0078125,-0.0078125,0.0546875,0.0546875,-0.03125,0.03125,0.0078125,-0.0234375,0,0.03125,-0.0625,-0.015625,0.0859375,0.0390625,-0.0390625,-0.0234375,0.078125,0.09375,-0.03125,-0.015625,-0.046875,-0.0078125,-0.0703125,0,0.0390625,0.0234375,-0.03125,0.0078125,-0.0078125,-0.015625,-0.0390625,0.0078125,-0.015625,0,-0.0234375,0.0078125,0,0.015625,0,-0.015625,-0.0390625,0.03125,0.1015625,-0.0546875,0,-0.0234375,0,0.0078125,0,-0.0546875,0,-0.0546875,0.0703125,0.03125,0.03125,-0.0625,-0.0625,-0.015625,0.1015625,-0.03125,-0.03125,0.0078125,0.046875,-0.0390625,-0.0078125,0.0546875,0.0078125,-0.0078125,-0.0078125,0.015625,0.0078125,0.0234375,0,0.0078125,0.0078125,-0.0234375,0.0078125,0.0234375,0.0390625,-0.0390625,0.015625,0.0625,0.015625,0,-0.0234375,-0.0703125,0.0078125,0.0078125,-0.03125,-0.0078125,0.0234375,0.03125,-0.046875,0.0078125,-0.09375,-0.0078125,-0.0703125,-0.109375,0,0.0546875,-0.0234375,0.078125,-0.0078125,-0.109375,-0.046875,0,-0.015625,0.0078125,-0.0234375,0.0546875,0.0390625,0.0078125,0,0.03125,-0.0390625,-0.0234375,0.0390625,0.0546875,0.015625,-0.015625,0,-0.015625,0.0390625,-0.0078125,-0.0078125,0.0234375,-0.0078125,-0.046875,0.0234375,-0.015625,-0.0234375,0.015625,-0.0546875,-0.109375,-0.0859375,-0.0234375,0,0.046875,0.0859375,0.03125,-0.0390625,0.03125,0.0234375,0.015625,0.0078125,-0.0234375,-0.0390625,0.0078125,0,-0.0234375,-0.0703125,0.03125,-0.015625,-0.0234375,0.046875,-0.0078125,-0.078125,-0.078125,0.0234375,0.015625,-0.0078125,0.015625,0.0078125,0,0.0078125,0.03125,0.1484375,0.0234375,-0.015625,-0.03125,-0.0546875,-0.03125,-0.03125,0,0.0546875,-0.0546875,-0.015625,0.015625,-0.0703125,-0.0625,-0.0234375,0.0703125,-0.0703125,-0.0859375,0.0703125,0.046875,-0.0703125,-0.0859375,0.03125,0.0546875,-0.0703125,0.0625,0.0078125,-0.0390625,0.0546875,-0.0234375,-0.03125,-0.0625,-0.0078125,0.0390625,-0.0234375,0.0078125,0.0859375,0.0390625,-0.09375,-0.078125,-0.015625,0.015625,-0.078125,0.015625,0.0078125,0.0234375,0.015625,-0.015625,-0.0390625,0.0078125,0.03125,0.0546875,0.0625,0,-0.015625,-0.015625,0,-0.0078125,-0.015625,-0.0078125,-0.0078125,0,0.0546875,0.015625,0.0703125,0.0390625,-0.0625,0.0078125,-0.03125,-0.015625,0,0.0234375,0.0546875,0.0078125,0.03125,-0.0234375,0,-0.0234375,-0.015625,-0.015625,0,-0.046875,0.0078125,-0.046875,0.03125,-0.015625,0.015625,0.0078125,-0.015625,0.0078125,-0.0078125,-0.0078125,-0.0078125,-0.015625,0.0078125,-0.0078125,0.0078125,0.0078125,0.03125,-0.015625,0,-0.015625,-0.046875,0.015625,0.0078125,-0.03125,0,-0.0234375,-0.046875,-0.0859375,0.0625,0.0390625,-0.015625,0.03125,-0.0078125,0.046875,0.0234375,-0.015625,-0.0234375,-0.0703125,-0.0078125,-0.015625,-0.0546875,-0.0625,-0.015625,0.015625,0.015625,-0.015625,0.078125,0,0.0078125,0,0,0.015625,0.0234375,0.0390625,-0.0234375,-0.03125,0.015625,-0.03125,-0.0078125,-0.046875,-0.0234375,-0.0078125,-0.0234375,-0.0234375,0.0078125,-0.0078125,-0.0078125,0.015625,-0.0078125,0.0078125,0,0.0078125,-0.0078125,-0.015625,-0.0078125,-0.015625,-0.0234375,0.0078125,0.046875,0.0234375,0,0.03125,0.0390625,-0.046875,0.0078125,-0.015625,-0.015625,-0.0234375,0,-0.03125,-0.0078125,0.0625,0.0390625,-0.0078125,0.03125,-0.0390625,-0.015625,-0.015625,-0.03125,0.0234375,0.0078125,-0.0234375,-0.015625,0.0390625,0.0234375,-0.046875,-0.0078125,0,-0.0078125,0,-0.015625,0.015625,-0.015625,-0.015625,-0.0078125,0,-0.0234375,-0.015625,0.0078125,0,-0.015625,0,0.0078125,0.03125,0.0078125,0.03125,0.0078125,0.046875,0.03125,-0.03125,0.0234375,0.015625,0.0234375,0.0234375,-0.03125,-0.03125,0.03125,0.03125,-0.03125,0,-0.0546875,-0.0234375,-0.015625,0.0078125,-0.0078125,0,0.03125,0.0546875,-0.0234375,-0.03125,-0.015625,0.015625,-0.03125,-0.03125,0.0234375,0.03125,-0.015625,-0.0078125,-0.0078125,0.0234375,0.0078125,-0.0078125,0.0078125,0.0078125,-0.015625,0.0078125,-0.0078125,0.0078125,0.015625,0.015625,0.0078125,0.1015625,-0.03125,-0.0625,-0.0234375,-0.03125,0.0234375,0.03125,-0.03125,-0.0234375,0.0078125,0,-0.0390625,-0.015625,0.0078125,0.015625,0.0078125,0.0078125,-0.015625,0.0078125,0,0.015625,0,-0.0234375,-0.0546875,0.0078125,0,-0.015625,-0.0234375,-0.03125,-0.0078125,-0.0078125,-0.015625,0.0078125,-0.0078125,-0.0234375,-0.0390625,0.015625,0.046875,-0.0546875,0.046875,-0.0078125,-0.046875,-0.03125,-0.03125,-0.0234375,-0.03125,-0.015625,0.0703125,-0.015625,0.015625,-0.0234375,-0.015625,0.0390625,0.0390625,0.0703125,0.015625,0,-0.015625,-0.0390625,-0.0546875,0.0078125,-0.0078125,-0.0703125,0.015625,0,-0.0078125,0.0234375,0.015625,0.0078125,0.03125,0.0078125,0.03125,-0.0078125,-0.03125,-0.0234375,-0.0703125,0.0078125,0.0390625,0.0625,-0.09375,0.0546875,0.015625,-0.0078125,0.0390625,0.015625,0.078125,0.09375,0,0.0078125,-0.0078125,0.0078125,0.0234375,0,-0.015625,0.015625,-0.0078125,-0.0078125,0.0234375,-0.0234375,0.03125,0.0546875,-0.0390625,-0.03125,0.0078125,-0.015625,0,0.0078125,-0.015625,-0.015625,0.0078125,-0.0234375,-0.0234375,-0.03125,-0.0546875,0.0078125,0.0234375,-0.0078125,-0.0078125,0.0234375,-0.015625,0.0234375,-0.0390625,-0.0546875,0,0,0,0.015625,-0.015625,-0.015625,0,0,-0.0078125,0.0078125,-0.0546875,0.015625,-0.015625,0.015625,0,-0.0234375,-0.046875,-0.0625,0,0.0234375,0.0234375,-0.0234375,-0.0234375,-0.0078125,0.0703125,0.0078125,-0.0546875,0.046875,0.0625,0,0.0078125,-0.0859375,-0.0078125,-0.0078125,-0.0546875,-0.0390625,-0.0078125,0.0078125,-0.0625,0.0078125,0.0078125,0.0625,-0.0390625,0.0078125,0.0390625,0.015625,-0.0703125,0.0703125,0.015625,0,-0.0625,0.0078125,-0.0390625,-0.03125,0.0234375,-0.0078125,0.03125,-0.03125,0,-0.0078125,0,-0.015625,-0.03125,0,-0.015625,-0.015625,-0.0078125,0.015625,-0.0234375,0.0078125,0.015625,0,0.0078125,0.046875,-0.0390625,0.0078125,-0.015625,-0.0546875,-0.0234375,-0.015625,-0.046875,0.0078125,0.0078125,0.015625,0.015625,-0.078125,-0.0390625,0.0078125,0.0390625,0.1015625,0.0859375,-0.0859375,0.0234375,-0.0234375,-0.0234375,-0.03125,-0.0078125,-0.015625,0,0.0234375,-0.0078125,0.0078125,0,-0.015625,0,0,0,0.015625,-0.0078125,-0.0078125,0.015625,-0.015625,0,0.0625,-0.046875,-0.015625,-0.03125,-0.03125,0.03125,-0.0078125,-0.0078125,-0.0234375,-0.0703125,-0.046875,0,0,-0.0390625,0.140625,0.015625,0,-0.1171875,-0.078125,-0.046875,-0.0703125,-0.03125,0,-0.078125,-0.0234375,0.0390625,-0.078125,-0.09375,0,0.046875,-0.0390625,0.0078125,0,0.0078125,-0.03125,0.0625,0.0546875,-0.046875,0.015625,-0.0078125,0,-0.0390625,0,-0.0390625,-0.015625,0.0390625,-0.03125,0.0234375,0,0,0.15625,-0.0625,-0.046875,0,-0.1015625,-0.0234375,-0.0546875,-0.0546875,-0.0625,-0.03125,0,-0.0234375,-0.0390625,-0.0234375,-0.046875,0,-0.015625,-0.0078125,-0.0703125,-0.0546875,-0.015625,-0.015625,-0.015625,-0.046875,-0.0078125,-0.0078125,-0.0234375,0.078125,-0.0078125,-0.0078125,0.015625,0,-0.0078125,-0.0546875,-0.0390625,0.0234375,0.0078125,-0.0078125,-0.0234375,-0.03125,-0.0078125,0,-0.0390625,-0.0234375,0.0625,-0.0078125,-0.046875,0.015625,-0.03125,-0.046875,0.046875,-0.03125,-0.03125,0.078125,0.015625,-0.015625,-0.015625,0.03125,0.03125,-0.0390625,-0.03125,-0.1015625,0.0234375,0,0,-0.015625,0.0703125,-0.0078125,0,0.0546875,-0.0078125,0.0234375,-0.078125,0.0078125,0,0.078125,0.0078125,0.0078125,-0.015625,-0.046875,0.0234375,-0.0234375,-0.046875,-0.0703125,0.0078125,-0.0078125,-0.0390625,0,0.0546875,-0.0234375,0.0078125,0.0078125,-0.0078125,0.015625,-0.015625,0.015625,0.015625,0.0078125,0.0078125,0,-0.03125,0,-0.0625,-0.0234375,0.0390625,0.03125,0.015625,0,0.015625,-0.0234375,0,0,-0.0234375,-0.0078125,0.0078125,-0.0390625,-0.0546875,-0.0390625,0.09375,-0.0078125,0.015625,-0.0078125,-0.0234375,0.0390625,-0.0078125,0.0078125,0.0078125,0.0078125,0,0,0.0078125,0,0.0078125,0.015625,0,0.03125,-0.0390625,-0.015625,-0.0078125,-0.03125,0.0546875,0.03125,0,0.0703125,-0.046875,-0.046875,0.0859375,-0.0390625,-0.0390625,0.0390625,0.015625,-0.1015625,0.0234375,-0.046875,0.0625,-0.0078125,-0.0390625,-0.0546875,-0.109375,-0.0078125,0.0390625,-0.03125,0,0.03125,-0.0078125,-0.0078125,0.015625,0,0,0.015625,-0.046875,-0.015625,0.0546875,-0.0390625,-0.0390625,-0.046875,-0.046875,-0.0078125,0.0859375,0.0546875,0.0234375,0.0234375,0.03125,0.0234375,-0.015625,0.015625,0.03125,0.015625,-0.015625,0.0390625,0.015625,0.046875,-0.0234375,-0.03125,0.015625,0,-0.015625,-0.0078125,0,-0.0078125,0.03125,0.0078125,-0.0546875,-0.046875,0.0078125,-0.0390625,-0.0625,0,0,-0.140625,-0.0390625,-0.0546875,0.0234375,-0.03125,0.046875,-0.0234375,-0.0390625,-0.0078125,0.109375,0.015625,-0.046875,-0.0703125,0.015625,0.0546875,0.0390625,0.0078125,0.015625,0.0078125,-0.0078125,0.0078125,0,-0.0078125,0,-0.0078125,0.0625,0.015625,0.03125,0,0.015625,-0.015625,0.0234375,-0.0234375,-0.0234375,0.0078125,0.015625,-0.03125,-0.0078125,-0.0859375,0.046875,0.0078125,0.0234375,0.015625,-0.03125,-0.03125,-0.0078125,-0.0234375,-0.0703125,0.2421875,0.0234375,0.0390625,-0.1171875,-0.0234375,0,0.0078125,-0.0234375,-0.0625,-0.015625,-0.0234375,-0.0390625,0.0078125,0,0.0546875,0,-0.03125,-0.0078125,-0.1015625,0.015625,0.0703125,0.0234375,0,0,0.0078125,-0.0078125,-0.03125,-0.046875,0.0390625,0.078125,0.0078125,0.0390625,-0.03125,0.0234375,-0.0078125,-0.046875,0.046875,0.0078125,0.015625,-0.0546875,-0.0234375,0.03125,0,0,0.0625,-0.0234375,0.015625,-0.0078125,-0.0390625,-0.015625,-0.046875,-0.0078125,-0.015625,0.015625,-0.046875,-0.015625,0.078125,0.09375,0.03125,-0.015625,0.0234375,-0.0234375,-0.0234375,-0.0390625,0.0703125,0.0234375,0.0390625,-0.015625,0.03125,0.015625,-0.0625,-0.0234375,-0.03125,-0.0078125,0,0.046875,0,0.046875,-0.0390625,-0.0234375,0.015625,0.0703125,-0.0390625,-0.0546875,-0.0859375,-0.0234375,-0.0390625,-0.078125,-0.0625,-0.03125,0,-0.046875,0.015625,0.0234375,-0.0390625,0.078125,0.0859375,-0.0234375,-0.03125,0.09375,-0.0078125,0.03125,0.015625,0.03125,-0.0625,-0.0078125,-0.0234375,-0.0390625,-0.03125,-0.0234375,0.078125,0.0859375,0.0078125,0.0546875,-0.0390625,0.015625,0.015625,0,-0.0546875,-0.0078125,-0.0234375,-0.0078125,0,0,0,0,-0.0078125,-0.0078125,0.0078125,0.0078125,0.0234375,0.0703125,0.0546875,-0.03125,-0.046875,-0.015625,0.046875,0.0859375,0.0234375,-0.0234375,-0.0390625,-0.0078125,-0.015625,-0.0546875,0.109375,0.015625,0.046875,-0.0234375,0.0078125,0,0.0390625,0.0390625,-0.015625,0.0234375,-0.0078125,-0.078125,-0.03125,-0.0078125,-0.0078125,0,0.015625,-0.0078125,0.0078125,0.0078125,-0.0078125,-0.0078125,0,-0.046875,-0.078125,-0.0703125,0.0078125,-0.015625,0.0546875,0.0859375,-0.03125,0.0234375,-0.0390625,-0.046875,-0.015625,0.0078125,0.0078125,0.0234375,-0.046875,-0.015625,-0.0390625,-0.03125,-0.0390625,-0.015625,0.0078125,0.0546875,-0.046875,0.0078125,-0.03125,0,0,0.0390625,-0.03125,-0.09375,-0.0234375,0.0390625,0.046875,-0.015625,-0.0234375,-0.03125,-0.015625,0.015625,0.0390625,0.0078125,-0.0078125,0.0390625,-0.0078125,-0.03125,-0.0546875,0.0546875,0,-0.015625,0.0078125,-0.015625,-0.03125,0.0390625,0.03125,-0.015625,-0.0078125,0,0.03125,-0.03125,0,-0.0234375,0.0078125,0.015625,0.03125,-0.015625,-0.03125,-0.0078125,0.015625,0,-0.0625,-0.046875,0.0234375,-0.0234375,-0.0546875,0.0390625,0.03125,0.078125,-0.046875,-0.0078125,-0.0625,-0.0390625,0.0546875,0.015625,0.03125,-0.0078125,-0.046875,0.0234375,-0.0078125,-0.0390625,0.0078125,0.0078125,0,0,0,0,0.0234375,0,0,0.015625,-0.03125,0,-0.0078125,-0.03125,-0.015625,0.0546875,0.0234375,-0.0078125,0.0625,-0.1328125,0.03125,0.0390625,0.03125,0.0078125,0.015625,-0.03125,-0.03125,0.03125,-0.0078125,-0.0546875,0.046875,-0.0546875,0.0625,0,0.015625,0,0.078125,0.0234375,0.0078125,-0.03125,-0.0390625,-0.0703125,0.0078125,0.015625,-0.0390625,0.0234375,-0.0078125,0.0546875,-0.0234375,-0.0546875,0.03125,0.0625,-0.0546875,0.0234375,0.0234375,-0.03125,-0.0078125,0,-0.03125,-0.0078125,-0.03125,0.03125,0.0078125,0.0625,-0.0625,0.03125,0.0703125,-0.0625,-0.015625,0.09375,-0.0078125,0.0390625,-0.03125,0.0234375,0.0234375,-0.0390625,0.0078125,0,0.0390625,0.015625,0.046875,-0.03125,-0.0078125,0.109375,0.03125,0.0078125,0.046875,0.03125,-0.0078125,0.0234375,-0.03125,0.0234375,0.0390625,-0.0546875,0.046875,-0.015625,-0.0234375,-0.046875,0.015625,0.046875,0.0546875,-0.0234375,-0.0625,0.0078125,-0.046875,0.046875,-0.0546875,0,0.0078125,0,-0.0234375,-0.0078125,0.078125,0.0078125,0.0078125,-0.0546875,-0.0078125,0.0390625,-0.0546875,0.0078125,-0.046875,-0.0390625,-0.0546875,0.03125,0.0078125,0.0390625,-0.015625,0.03125,-0.046875,-0.0234375,0.0390625,-0.0390625,-0.03125,0.0078125,0.0078125,0.1171875,-0.09375,-0.015625,0.0625,-0.046875,-0.0234375,0.0234375,0,0.015625,0.03125,-0.09375,-0.0546875,-0.046875,0.0078125,-0.0078125,0.03125,-0.015625,-0.0390625,0.0078125,0.0078125,0,-0.015625,0,0,0,0.015625,0,0.0234375,0,0,0,0.0078125,-0.078125,-0.0625,0.0078125,-0.0234375,-0.03125,0.015625,0,0,-0.0625,-0.015625,0.0078125,0,0.0078125,0.0625,0.0390625,0.0234375,0.046875,0.03125,-0.015625,-0.0234375,-0.046875,-0.0078125,0.015625,-0.015625,0.0078125,0,0,0.0078125,0.0078125,-0.0078125,0,-0.015625,-0.0078125,0.015625,-0.0078125,-0.125,0.078125,0.0078125,0.0703125,-0.09375,0.015625,0.0546875,-0.015625,0.0703125,0.046875,0,-0.046875,0.03125,0.0546875,0.015625,0.0390625,0.0390625,-0.0234375,0,-0.09375,0.0234375,0,0.015625,-0.0234375,0,0,-0.015625,0.046875,-0.09375,0,-0.015625,0.015625,-0.03125,0.03125,-0.0078125,0.046875,-0.0234375,0.046875,0.0625,-0.0078125,-0.03125,0.03125,-0.015625,-0.0234375,-0.0546875,0.0390625,-0.0078125,-0.03125,-0.015625,0.0234375,-0.0078125,0.0390625,-0.015625,-0.015625,-0.015625,-0.0078125,-0.03125,0.015625,0.0390625,0.0625,0.0234375,-0.0234375,-0.0390625,-0.0390625,-0.03125,0.0234375,0.03125,-0.0078125,-0.078125,-0.0625,0,-0.0234375,-0.0390625,0.0078125,0.0703125,0.0234375,-0.015625,-0.015625,-0.0078125,0,0.109375,-0.046875,-0.046875,-0.046875,-0.015625,-0.0703125,0,-0.0078125,0,0.015625,0,-0.015625,0,-0.015625,-0.0078125,0,-0.015625,-0.015625,-0.0390625,0.0078125,-0.015625,0,-0.015625,-0.0625,-0.0078125,-0.0234375,-0.0078125,-0.0234375,0.078125,-0.0078125,0.015625,-0.0390625,0.0078125,-0.0234375,0.046875,0.0078125,-0.0078125,0,-0.0234375,-0.0078125,-0.015625,-0.0234375,0.0234375,-0.0703125,-0.015625,-0.0078125,0.03125,0.0078125,0.015625,0,-0.015625,0.0390625,-0.03125,-0.0390625,-0.0546875,0,-0.0390625,0.0703125,-0.0625,0.015625,0.09375,-0.0078125,0.015625,-0.015625,-0.0390625,-0.0390625,-0.0078125,-0.046875,0.015625,-0.0390625,0.046875,0.015625,-0.0078125,-0.0546875,0.0859375,-0.0703125,0.0078125,0.0078125,-0.0078125,0,-0.0234375,-0.046875,0.0390625,-0.0625,0.0234375,0.0546875,-0.015625,-0.015625,-0.0078125,0.0078125,-0.03125,0.0234375,-0.0078125,-0.0546875,0.125,0.1015625,0.046875,0.078125,-0.046875,-0.0078125,-0.0546875,-0.0546875,-0.03125,0.015625,0.0625,-0.0390625,0.0078125,-0.0078125,0.1015625,-0.125,-0.0390625,0.0234375,0.0078125,-0.015625,-0.0078125,-0.0234375,0.03125,0.0859375,0.0546875,0.0546875,-0.03125,-0.0234375,-0.046875,0.015625,0.0390625,0.03125,-0.015625,-0.0234375,-0.03125,-0.015625,0.1171875,0.015625,0.03125,0.0703125,0.0625,0.0234375,-0.03125,-0.0234375,-0.046875,-0.0234375,-0.0390625,0.0078125,0.0078125,0.0234375,-0.0078125,-0.015625,0.0625,0,-0.0234375,-0.0078125,-0.0078125,0.0234375,0.0078125,0.0234375,-0.0546875,0.140625,0,-0.046875,0.0078125,-0.0078125,0.015625,-0.0078125,0,0.03125,0,-0.0078125,0.0234375,0,-0.015625,0,0.078125,-0.1015625,0.015625,0.0390625,-0.0703125,-0.0078125,-0.03125,-0.0546875,-0.0546875,0.015625,0,-0.0390625,0.0234375,-0.0234375,0.015625,0,-0.0546875,0,-0.0390625,-0.046875,0.03125,0.0078125,0,-0.0625,0.03125,0.015625,-0.015625,-0.0078125,-0.015625,-0.0078125,0,0.0078125,0,0.0078125,0.1171875,0.0703125,0.0859375,-0.03125,-0.15625,0.0546875,0.0234375,-0.0390625,0,-0.03125,-0.0390625,-0.03125,0.1015625,0.015625,-0.0390625,-0.0234375,-0.0703125,0.046875,-0.03125,0.1328125,-0.0390625,-0.0390625,0.0859375,-0.140625,-0.046875,-0.046875,-0.078125,0.03125,-0.03125,0.0078125,-0.0078125,-0.03125,0,0.0234375,-0.0546875,-0.0234375,0.046875,0.125,-0.0078125,-0.046875,-0.015625,0,-0.015625,0,0,0.0078125,-0.03125,0.03125,0.046875,-0.03125,0,0.03125,-0.0078125,0.03125,0,-0.0546875,0,0,0,-0.046875,0,-0.0078125,0.0234375,-0.015625,-0.0078125,-0.0546875,-0.03125,0.0234375,-0.0234375,0.0234375,0.03125,-0.0078125,-0.015625,0.0546875,0.015625,-0.0703125,0.046875,0.0234375,-0.078125,-0.1015625,0.0078125,-0.0703125,0.0234375,0.0703125,-0.0625,0.0625,-0.0078125,-0.0234375,0.015625,-0.046875,-0.0078125,0.0078125,0.0078125,-0.015625,-0.0078125,0.015625,-0.0078125,0,-0.015625,-0.0234375,-0.046875,0.0234375,0,-0.0390625,0,0,-0.046875,0.046875,0.0390625,-0.1171875,-0.046875,0.015625,-0.015625,-0.0078125,-0.0703125,-0.015625,0.015625,-0.015625,0.0859375,-0.0546875,-0.0078125,0.0390625,0.015625,0.015625,-0.03125,0.0234375,-0.0625,0.1015625,0.0078125,-0.0390625,-0.0546875,0,-0.0078125,-0.046875,0.0859375,-0.0625,-0.0625,-0.0078125,-0.0546875,-0.0625,-0.0078125,-0.0390625,-0.0078125,-0.046875,0.015625,-0.03125,0.078125,0.078125,-0.0078125,-0.0078125,-0.0234375,-0.015625,-0.078125,-0.140625,0.046875,-0.015625,-0.046875,0.0859375,-0.078125,-0.015625,-0.03125,-0.0078125,-0.0703125,0.0390625,-0.046875,-0.0546875,0.015625,-0.125,-0.015625,0.09375,0.015625,-0.0625,0.0390625,-0.0546875,-0.03125,-0.0078125,-0.03125,-0.0625,0.0390625,-0.0234375,0.0078125,-0.0625,-0.0625,0.0234375,0.015625,0.0234375,-0.0390625,-0.0390625,-0.03125,0.0078125,0.03125,0.046875,-0.0390625,0,0,-0.03125,0.0546875,-0.0546875,-0.0390625,0.015625,0.09375,-0.046875,-0.0546875,-0.1171875,0.03125,0.1015625,0.109375,-0.0234375,0.0625,0.046875,-0.0546875,-0.0390625,-0.0078125,-0.03125,0.015625,-0.046875,-0.0234375,-0.0625,0.0625,-0.03125,0.0078125,0,0.0234375,0.0234375,0.109375,0.15625,-0.0546875,0.0234375,0.0390625,-0.03125,0.0390625,-0.0234375,0.0078125,0,0.046875,-0.0390625,-0.0390625,-0.03125,0.0546875,-0.046875,0.109375,0.0078125,0.0625,0.0078125,-0.0078125,0.015625,-0.0078125,0.0078125,-0.015625,0,0.0078125,0.015625,0.0078125,0.0625,0.0078125,-0.0859375,0,-0.03125,0.0546875,-0.046875,-0.0078125,-0.0390625,-0.0703125,0.0078125,-0.0234375,-0.015625,-0.0234375,0.0703125,-0.0625,-0.0703125,-0.0078125,-0.0078125,-0.046875,0.0625,-0.0234375,-0.046875,-0.0234375,0.03125,-0.015625,0.0078125,-0.0078125,-0.015625,-0.0078125,0,0.0078125,-0.0078125,-0.0078125,-0.0078125,0,0.0546875,0.015625,-0.0234375,-0.046875,-0.078125,-0.0546875,-0.125,-0.0234375,0.015625,0.09375,-0.078125,0,-0.015625,-0.0390625,0,0.015625,0,-0.1015625,-0.0625,-0.0625,0.0078125,0,0,0.0625,-0.0078125,-0.0390625,0.0234375,-0.03125,0.0390625,0.0234375,-0.0234375,-0.0859375,0.015625,0.046875,-0.0234375,-0.0390625,0.046875,-0.0078125,-0.0703125,0.015625,0.0234375,0.0234375,-0.0546875,0.0234375,-0.078125,-0.046875,-0.03125,0.0078125,0,0.0078125,-0.0234375,0.0078125,0.015625,-0.0546875,0,0.0078125,-0.0234375,-0.0234375,0.03125,0.015625,-0.015625,0,-0.0234375,-0.0234375,0,-0.0546875,-0.015625,-0.015625,-0.0625,-0.03125,-0.046875,0.0078125,0,-0.03125,0.046875,0.015625,0.0546875,0.171875,-0.0703125,0.015625,0.015625,0.0625,0,-0.0390625,-0.0234375,-0.0234375,0.1328125,0.03125,-0.015625,-0.0078125,-0.0078125,0.0078125,0.015625,-0.015625,0.0078125,0,-0.03125,0,0,-0.015625,0,-0.0234375,0.03125,-0.046875,0,-0.0703125,0.0078125,-0.0703125,-0.046875,-0.0703125,-0.03125,0.0625,-0.0078125,-0.0625,0.0078125,-0.046875,-0.046875,0.0390625,-0.03125,-0.0546875,-0.03125,-0.0078125,0.0390625,-0.0625,0.0703125,0.0078125,-0.015625,-0.015625,0.046875,-0.0234375,-0.0703125,-0.03125,-0.0234375,-0.046875,-0.03125,-0.0390625,0.0234375,-0.078125,0.03125,0.0078125,0.0625,0.171875,0.0078125,-0.0390625,0.0703125,-0.03125,-0.03125,0.1484375,-0.0390625,-0.0546875,-0.03125,0.015625,0.03125,-0.078125,-0.046875,-0.1015625,0.1015625,0.03125,-0.0703125,-0.015625,-0.0625,0.0234375,-0.0234375,0.03125,-0.015625,-0.015625,0.0078125,-0.0234375,-0.0390625,0.0078125,-0.0625,-0.046875,-0.046875,0.015625,-0.0625,0,-0.0625,-0.015625,-0.0625,-0.078125,-0.0390625,-0.0234375,0.015625,0.046875,0.03125,-0.015625,-0.0078125,-0.078125,0.0234375,-0.0390625,-0.03125,0.0078125,-0.09375,0.0625,-0.0546875,-0.046875,-0.015625,-0.046875,0.03125,-0.0625,0,0.03125,0.0234375,0.09375,0.03125,-0.046875,-0.046875,0.03125,-0.0234375,-0.046875,-0.1015625,0,-0.046875,0,0.0078125,-0.0546875,0.1796875,-0.03125,-0.0859375,0.09375,0,0,-0.109375,-0.0546875,-0.0234375,-0.0703125,-0.0078125,-0.0703125,0.0625,-0.015625,-0.015625,0,-0.03125,0.0234375,-0.046875,-0.0078125,-0.0546875,0.0546875,0.015625,-0.0234375,-0.0390625,0.0390625,0.0078125,0,0.0078125,0.015625,-0.015625,-0.0078125,0,0,-0.0078125,0.03125,-0.046875,-0.0390625,0.015625,-0.0078125,0.03125,-0.0078125,-0.015625,-0.015625,0,0.0078125,-0.03125,0,-0.0078125,0.0234375,0,-0.0078125,-0.0546875,0.03125,0.03125,-0.0390625,-0.0546875,0.015625,0.078125,-0.0234375,0,0.015625,0,-0.0078125,-0.0078125,0.0078125,0.0078125,0.0078125,0.0078125,-0.0078125,0.015625,0.03125,0,0,0.046875,-0.0078125,-0.015625,0.015625,-0.0546875,-0.0234375,-0.0078125,-0.0390625,0,-0.0234375,0.0390625,-0.03125,-0.0625,-0.03125,-0.03125,-0.0390625,-0.015625,0.0078125,-0.0859375,0,0.0703125,-0.015625,0.015625,-0.0546875,0.03125,-0.03125,0.015625,-0.0390625,-0.0390625,-0.0078125,0,-0.0078125,-0.0078125,-0.015625,-0.0625,-0.0546875,0.0390625,-0.0390625,-0.015625,0.0234375,0.0078125,0.03125,0,-0.0078125,-0.015625,-0.0078125,-0.0234375,0.015625,-0.015625,-0.0078125,-0.0078125,0.0078125,-0.0078125,-0.0078125,-0.0078125,-0.0078125,-0.015625,-0.015625,-0.03125,0,-0.046875,-0.0078125,-0.03125,-0.03125,-0.0390625,0.046875,-0.0078125,0.0078125,-0.015625,0.0390625,0.0078125,-0.046875,0.0390625,0,-0.015625,0.015625,0.0234375,0.0234375,0.015625,-0.0078125,0.078125,-0.0234375,0.015625,0.0234375,0.0234375,0.0078125,0,0.015625,0.015625,0,-0.0078125,0.015625,0.03125,0,-0.0078125,-0.0078125,-0.03125,0,-0.0390625,0,0.0234375,-0.0390625,0.0234375,0.015625,0.0390625,0.0078125,0.0234375,0.015625,0.046875,-0.0234375,-0.0234375,-0.046875,-0.0546875,-0.03125,0.046875,-0.0078125,-0.015625,0.0234375,0.015625,0.03125,0.015625,-0.0234375,-0.0546875,0.046875,0,-0.0078125,0.015625,0.03125,-0.0625,-0.03125,-0.03125,-0.0234375,0.0078125,-0.0078125,-0.0078125,-0.0546875,-0.0390625,0.0234375,-0.015625,-0.015625,0,0.078125,0.015625,-0.0234375,0.0546875,-0.015625,0,0.015625,0.015625,-0.03125,-0.03125,0,0.046875,0.078125,0.0078125,-0.0625,-0.0234375,-0.0078125,-0.0546875,-0.03125,0.0234375,-0.09375,-0.0234375,0.046875,0.0390625,-0.0078125,0.0859375,0.0625,0,0,-0.0234375,-0.0390625,0,0.03125,-0.015625,0.015625,0.046875,0.03125,0.0390625,-0.015625,0.015625,0.1015625,0.0390625,-0.03125,-0.0390625,-0.0234375,-0.1015625,-0.046875,0.1015625,-0.0234375,-0.0078125,0.0390625,0.0234375,-0.03125,-0.0546875,0.0078125,-0.078125,-0.046875,0.046875,0.078125,-0.0625,-0.03125,-0.046875,0.015625,-0.03125,-0.1015625,-0.0390625,0.0078125,-0.0703125,0.0234375,-0.015625,-0.046875,0,0.015625,0.03125,-0.046875,0.03125,-0.0234375,-0.0390625,0.0078125,0,-0.0078125,-0.078125,-0.046875,0,-0.03125,-0.03125,0.0390625,0.0078125,-0.0078125,-0.015625,0.015625,0,-0.046875,0.0625,0.0546875,-0.03125,-0.0390625,-0.0078125,0,-0.0078125,0.015625,0.015625,0,0.015625,0,-0.015625,-0.015625,0,0.0390625,-0.0234375,0,0.0546875,-0.0234375,0.0078125,-0.0234375,0.015625,0.015625,0.046875,0.015625,0.0078125,0.015625,-0.015625,-0.0546875,-0.0234375,-0.015625,0.078125,-0.03125,0.03125,0.0390625,-0.0078125,0.046875,-0.0078125,-0.015625,-0.0234375,0,0.0078125,-0.0078125,0.0078125,0,-0.0078125,-0.0078125,-0.0078125,-0.0078125,0.0078125,-0.015625,0,-0.03125,0,-0.046875,0.015625,-0.03125,0,0.0546875,0,-0.03125,-0.0625,0.109375,-0.015625,-0.0078125,-0.0625,0.0078125,0.0234375,0.03125,-0.015625,0.015625,-0.0078125,-0.0390625,0.015625,-0.0625,-0.0078125,0.03125,0,-0.0234375,-0.0078125,0,-0.046875,0.0625,0.0234375,0.03125,0.0078125,0.0078125,0.0078125,-0.03125,-0.03125,0.0078125,0.046875,-0.0390625,-0.015625,0.015625,-0.0078125,-0.015625,-0.015625,-0.046875,-0.046875,0.015625,0,-0.0234375,-0.03125,0.0078125,0,-0.0234375,0.03125,0.0078125,-0.0390625,0,-0.015625,0,0,0.015625,-0.015625,0.015625,-0.0078125,0.0078125,-0.0234375,-0.03125,-0.0078125,-0.0546875,-0.03125,0.0234375,-0.03125,-0.0078125,0.0703125,-0.015625,-0.03125,0.015625,-0.046875,-0.0390625,0.0703125,-0.03125,-0.03125,0.046875,-0.0234375,-0.03125,-0.0625,0.0078125,-0.015625,0.0078125,0,-0.0078125,0,0.0078125,0,0,-0.015625,0.0078125,0.03125,-0.03125,-0.015625,-0.03125,0,0.0234375,0.03125,-0.046875,-0.0234375,0.0625,0.0625,-0.015625,-0.0546875,0.03125,-0.015625,-0.0078125,-0.015625,-0.046875,-0.015625,0.0234375,0.0546875,0.0390625,-0.0078125,-0.0078125,0.09375,-0.0234375,0,0.078125,0.015625,-0.0234375,-0.0703125,0,-0.0390625,-0.0546875,-0.0234375,0.015625,0.0234375,0.015625,0.046875,0.0390625,-0.0625,-0.046875,-0.015625,0.0390625,0,-0.046875,0.046875,0.0234375,-0.03125,-0.046875,-0.0234375,-0.0234375,-0.03125,-0.0390625,0.0546875,0.03125,-0.0546875,-0.0859375,0.03125,0.0234375,-0.0625,0.03125,0.0234375,-0.03125,-0.0078125,0.0078125,0,-0.0078125,0.015625,0.015625,0.0234375,0.015625,-0.0078125,-0.0078125,-0.0078125,0.046875,-0.03125,-0.0546875,-0.0390625,0.0078125,0.0078125,0.03125,-0.03125,0.03125,0.0078125,-0.0234375,-0.0390625,0.0078125,-0.03125,-0.0703125,0.0390625,-0.046875,-0.03125,0.0703125,-0.015625,-0.046875,-0.03125,0,-0.015625,0.03125,0.015625,0,-0.046875,0.0625,0,0.03125,0.0234375,-0.015625,0.0390625,0.0546875,-0.046875,-0.0234375,-0.0234375,-0.015625,-0.0078125,0.0078125,0.0234375,-0.015625,0.0546875,0.0078125,-0.0625,0,0.015625,0.0078125,0.015625,0.046875,0.0546875,0.03125,-0.0234375,-0.0390625,-0.0234375,0,0,-0.0390625,0.015625,-0.0234375,-0.0078125,0.0078125,-0.0546875,0.0078125,0,-0.03125,0,-0.015625,0,-0.0078125,0,0.0234375,0.015625,-0.0078125,0,0.0859375,0.015625,-0.0078125,0.0234375,0,-0.0078125,0.03125,0.0234375,-0.0078125,0.078125,0.015625,-0.03125,0.046875,0.015625,-0.0078125,-0.0078125,0.0390625,0.0078125,-0.03125,-0.03125,-0.015625,-0.015625,0.046875,-0.0078125,0,-0.0546875,-0.0234375,-0.0078125,-0.0078125,0,0.0078125,0.0078125,0.0078125,0.0078125,0.0078125,-0.0078125,0.015625,0.1015625,0.015625,-0.046875,-0.0546875,-0.0078125,-0.0546875,0.0078125,-0.0390625,0.0546875,-0.0546875,0.03125,-0.0390625,0.046875,0,-0.0078125,-0.03125,-0.0546875,-0.03125,-0.0234375,0.0234375,-0.0625,0.1328125,0.0078125,-0.015625,0.046875,-0.0078125,0,0.015625,-0.0078125,0.03125,-0.015625,0,0,-0.0390625,-0.015625,0.0234375,-0.0078125,0.03125,-0.0859375,0.0390625,0.078125,-0.015625,-0.0234375,-0.0078125,0,-0.0390625,-0.03125,0.0390625,-0.015625,-0.0390625,0,-0.0078125,0.046875,0.03125,0.0390625,0.03125,0,0,0.03125,-0.0234375,-0.0078125,0.0390625,0.0234375,-0.0078125,-0.03125,0.015625,-0.0625,-0.0234375,-0.0078125,0.0078125,0,-0.03125,-0.0625,0.015625,-0.0078125,-0.0078125,-0.0546875,0.0078125,0.0078125,0.046875,-0.0625,-0.0625,0.0234375,0,0.0859375,0.03125,0,-0.0390625,-0.046875,0.0078125,0,0,-0.0078125,-0.015625,0.0078125,-0.0078125,0,0,0.078125,-0.015625,-0.03125,-0.0234375,-0.0234375,-0.0234375,0.0078125,-0.0078125,-0.015625,-0.0234375,0,-0.0390625,-0.015625,0,-0.015625,0.0390625,0.0703125,-0.03125,-0.0703125,-0.046875,0.125,0.0078125,-0.046875,-0.1015625,0.0546875,-0.0546875,-0.0078125,0.046875,0,-0.0390625,-0.0390625,-0.0546875,0.0546875,-0.03125,0.015625,-0.03125,0.015625,0.0625,0.0078125,0.0625,-0.0703125,-0.015625,0.015625,-0.0703125,-0.0078125,0,0.0234375,-0.0234375,-0.015625,0.0390625,-0.0390625,0.015625,0.0390625,0,0.03125,-0.0390625,0.046875,0.015625,0,-0.046875,-0.03125,0.046875,-0.0078125,-0.0078125,-0.046875,-0.0078125,-0.03125,-0.0234375,-0.0234375,0.0390625,0.0546875,0.0703125,-0.015625,-0.0078125,-0.0390625,-0.03125,-0.015625,0.03125,0.015625,0.03125,-0.0078125,0.046875,-0.0234375,0.0390625,0.03125,-0.0546875,-0.0234375,0.015625,-0.0546875,0.0078125,0.0390625,-0.078125,-0.0390625,0,-0.03125,-0.0703125,-0.0078125,0.0234375,0,0.015625,0.03125,-0.0390625,-0.0390625,-0.015625,0.0078125,-0.03125,0.0234375,0.0078125,0.09375,0.03125,0,0,-0.0625,0.03125,-0.03125,-0.0078125,0.0078125,0.0390625,0,0.03125,-0.0078125,-0.046875,0.0625,0.0234375,0,-0.0234375,-0.0234375,-0.0234375,0,-0.0546875,0,-0.0390625,-0.046875,0.0234375,0.015625,0,-0.0625,-0.0078125,-0.0078125,0.015625,0.0234375,0.0234375,-0.0390625,-0.015625,-0.015625,-0.0078125,0,-0.0078125,0,0.015625,0,0.0078125,-0.0078125,0.0078125,0.0625,0.0078125,0.0546875,-0.015625,-0.015625,0.015625,-0.0390625,0.0078125,0.0234375,-0.0703125,0.03125,0.0234375,0.1015625,-0.046875,0.0078125,-0.015625,-0.0546875,0.078125,0.0703125,-0.0234375,-0.0703125,-0.0703125,0.0078125,-0.0546875,-0.0078125,-0.0078125,0.015625,0,0,0.0078125,-0.0078125,0,-0.0078125,0.0078125,0,-0.0078125,-0.015625,0.046875,0.0390625,-0.0234375,-0.0546875,0.0078125,0,-0.015625,-0.0625,-0.015625,-0.0625,0.0390625,0.046875,0.0390625,0.09375,-0.03125,0.015625,-0.0234375,-0.0546875,0.015625,0.03125,0.0234375,0.015625,-0.03125,-0.0625,-0.0234375,-0.0078125,-0.0078125,0.0078125,-0.0078125,-0.0390625,-0.0078125,0.0390625,0,0.0078125,0.0078125,0.0078125,0.0078125,-0.03125,0,0.015625,-0.0703125,-0.0390625,0.0078125,-0.015625,-0.0078125,-0.03125,-0.0078125,-0.015625,-0.0078125,-0.015625,-0.015625,-0.0078125,-0.0234375,0,-0.0390625,0.0078125,-0.015625,-0.015625,0,-0.0078125,0.015625,0.0234375,-0.0390625,-0.03125,0.0078125,-0.03125,0,-0.0078125,-0.0078125,-0.03125,-0.0078125,-0.0546875,0.0390625,0,0,0.0078125,0.0859375,-0.0078125,-0.0234375,0.0546875,0.015625,-0.0078125,-0.046875,0.0078125,0.0546875,-0.0390625,-0.015625,-0.0234375,0.015625,0.015625,0.0078125,0,-0.0078125,0,-0.0078125,-0.015625,-0.0078125,0.03125,0,0.03125,-0.0078125,0.0078125,-0.015625,0.0234375,-0.03125,0.0546875,-0.03125,-0.0078125,-0.046875,-0.03125,0.046875,-0.0625,-0.015625,0.015625,-0.0234375,-0.046875,-0.0078125,0.0234375,0.03125,-0.0625,-0.0703125,0.0078125,-0.015625,0.0234375,0,-0.0390625,-0.0234375,-0.0078125,0,-0.0078125,-0.015625,-0.0234375,-0.03125,0,0.1015625,-0.03125,-0.046875,-0.0859375,-0.015625,-0.0078125,0.0234375,0.0390625,0.0078125,-0.015625,0.0078125,-0.0078125,0.0625,-0.046875,-0.0234375,0.046875,-0.0390625,-0.0234375,0.0546875,-0.0078125,-0.046875,-0.03125,-0.0390625,-0.0078125,0,-0.078125,0.0859375,0,-0.0234375,-0.0390625,-0.015625,-0.0625,-0.0546875,0,0.03125,-0.0234375,0,-0.015625,-0.03125,0.046875,0.015625,-0.046875,0.078125,0.0546875,-0.015625,-0.0078125,-0.0390625,0.015625,0.0859375,-0.0234375,-0.015625,-0.0625,0.0234375,-0.03125,0.0078125,0.0703125,-0.0078125,-0.09375,0.0390625,-0.0078125,-0.0625,0,0.0625,-0.0234375,0.046875,0.0546875,-0.0234375,-0.0078125,-0.0625,0.015625,-0.0078125,-0.046875,0.03125,-0.0078125,0.0078125,0.0390625,-0.015625,-0.015625,-0.0390625,-0.015625,-0.046875,-0.015625,0.03125,-0.0078125,0.03125,-0.03125,0.03125,0.0078125,-0.0234375,-0.0234375,0.0234375,-0.0078125,-0.0390625,-0.0078125,-0.03125,-0.0078125,0.078125,-0.015625,-0.0703125,-0.0234375,-0.0078125,-0.046875,0.015625,0.015625,-0.0234375,-0.0078125,0.0234375,0.015625,0,0.0078125,0.015625,-0.0078125,-0.015625,-0.0078125,0.0078125,0.015625,0.0546875,-0.015625,0.015625,0.015625,0.015625,0.03125,-0.015625,-0.015625,-0.03125,0.0078125,0.046875,0.046875,-0.0390625,-0.0078125,-0.015625,-0.015625,0.015625,-0.015625,0.0078125,0.0078125,-0.046875,0.046875,-0.015625,-0.0078125,0,-0.015625,-0.0234375,0.0078125,0,-0.0078125,0.0078125,0,0.0078125,0,-0.0078125,-0.015625,-0.03125,0.015625,-0.015625,0.046875,0.046875,-0.03125,-0.015625,-0.0234375,-0.015625,0.125,-0.03125,-0.015625,-0.078125,-0.03125,-0.03125,-0.0078125,-0.0234375,0.0078125,-0.0234375,0.0078125,0.03125,-0.0625,-0.0078125,-0.0546875,-0.0078125,-0.03125,-0.015625,0.015625,-0.0078125,0,0.0078125,0.015625,0,-0.0078125,-0.0234375,0.015625,-0.0078125,0.0078125,-0.0078125,0.0234375,-0.0234375,-0.03125,-0.03125,-0.015625,0.015625,0.0078125,0.0234375,-0.0078125,0.0390625,-0.0390625,-0.0078125,0.0078125,-0.0234375,-0.0078125,0.0078125,-0.015625,-0.015625,-0.0078125,0,0,0.0078125,-0.0078125,0.015625,0.0078125,0.015625,0,-0.078125,-0.015625,0,0.015625,0,0,0.125,-0.046875,-0.03125,-0.1015625,-0.046875,-0.03125,-0.0078125,0,0,-0.0859375,0.0546875,-0.0546875,-0.03125,-0.0078125,0,-0.0078125,0.0078125,0.0390625,-0.0234375,-0.015625,0.015625,0,-0.0078125,-0.0078125,0.0078125,0,-0.0078125,-0.0234375,0.0078125,-0.0078125,-0.015625,0.03125,0.03125,-0.015625,0,-0.0078125,0.0625,-0.078125,0.015625,0.0078125,0.015625,0.0078125,-0.03125,0.0234375,0.03125,0.2890625,0.0703125,-0.0390625,-0.1875,-0.046875,-0.0625,-0.0390625,-0.0078125,-0.0078125,0.03125,-0.0390625,-0.015625,-0.03125,0.015625,0.0234375,-0.03125,-0.0078125,0.0078125,-0.0390625,-0.0234375,-0.015625,0.03125,-0.0078125,0.0390625,-0.0390625,-0.0625,0,-0.015625,-0.0625,0,0.0078125,0.046875,0.0703125,-0.0078125,0,0.0078125,0.1015625,-0.015625,0.0390625,-0.03125,-0.0859375,0,-0.015625,-0.0078125,0,0.0390625,0.0234375,-0.0078125,0.015625,-0.0859375,-0.0234375,-0.0234375,-0.0390625,0.015625,-0.0078125,-0.0390625,0.0234375,0.03125,0.03125,0.046875,0.015625,0,-0.0234375,-0.0078125,0.0078125,-0.03125,-0.0546875,-0.015625,-0.0546875,0.015625,-0.0078125,-0.015625,0.0703125,-0.0078125,-0.03125,-0.046875,-0.0390625,0,-0.015625,0.03125,-0.03125,0.1015625,-0.0390625,0.0078125,-0.0234375,-0.0625,-0.0078125,-0.0234375,-0.015625,0.03125,0.03125,0.03125,0.0234375,0.015625,0.015625,0.0234375,-0.0234375,-0.046875,-0.015625,0.015625,-0.0625,-0.0234375,0.03125,-0.0234375,0.0546875,-0.0234375,0.015625,0.015625,-0.0234375,-0.046875,-0.015625,-0.015625,-0.046875,0.03125,-0.0234375,-0.0078125,0.0234375,-0.015625,-0.0390625,0.0078125,0.125,-0.0078125,-0.0234375,-0.0234375,0.03125,-0.0078125,-0.015625,-0.0078125,0.0078125,0.015625,0,0,0.015625,0,0.0078125,0,0.0234375,-0.0078125,0.03125,-0.0859375,-0.046875,-0.0234375,-0.0078125,-0.0234375,-0.03125,-0.015625,0.0390625,-0.0234375,0.0625,0.03125,0,0.0078125,-0.015625,-0.0390625,0.046875,-0.0078125,-0.0390625,0,0.015625,0.1171875,0.0390625,-0.015625,0,0.0078125,-0.0078125,0,-0.0078125,0,-0.0078125,-0.0078125,0.0078125,-0.015625,0,-0.03125,-0.0234375,-0.0703125,-0.015625,0,-0.0625,-0.0390625,0.0234375,0.0234375,-0.0078125,0.0078125,0.0625,-0.0078125,0.0234375,0.0234375,-0.015625,-0.09375,-0.046875,0.078125,0.03125,-0.0390625,0.015625,0.0546875,-0.015625,-0.0234375,0.0625,-0.0078125,-0.0234375,0.046875,0.0078125,-0.0546875,-0.0546875,0.015625,-0.0234375,0.015625,-0.0234375,-0.0390625,0.0625,0,-0.015625,0.0390625,-0.0078125,-0.015625,0.03125,-0.03125,-0.0234375,0.046875,0.0234375,0.0390625,-0.03125,-0.015625,0.0078125,-0.03125,0.0234375,-0.0078125,-0.015625,-0.0078125,0.015625,0.0078125,0.0234375,0.015625,0.0078125,0.0078125,0,0.0234375,-0.015625,0.03125,0.015625,-0.0703125,-0.0234375,-0.0234375,-0.0703125,-0.0390625,0,0.0546875,-0.046875,0.0078125,0.0078125,-0.015625,-0.03125,-0.03125,-0.03125,-0.125,-0.0078125,0.0078125,0.0703125,0.09375,-0.0078125,-0.0078125,-0.0078125,-0.0078125,-0.015625,0,0.0078125,0.03125,0.03125,-0.0078125,0.03125,0.0390625,0,0.0078125,-0.046875,0,0.0078125,0.0234375,-0.0078125,0,-0.0078125,-0.0234375,-0.0390625,0.0546875,-0.015625,0.015625,0.0546875,-0.015625,-0.03125,-0.0390625,-0.0234375,-0.1015625,-0.046875,-0.0390625,0.0546875,0.0078125,-0.0078125,0.0078125,-0.078125,-0.0390625,-0.0390625,-0.0390625,0.0078125,0.1015625,0.0859375,-0.0234375,0.03125,0.0703125,-0.0390625,-0.109375,0,-0.015625,-0.0234375,0.0390625,-0.046875,-0.0703125,0.03125,0.0234375,0.046875,-0.0078125,-0.03125,0.015625,-0.015625,0,0.015625,-0.0078125,-0.015625,-0.015625,-0.015625,-0.0234375,0.0390625,-0.1015625,-0.0234375,0.03125,-0.03125,0,-0.046875,-0.03125,-0.015625,-0.0234375,-0.0078125,-0.0234375,0.0390625,-0.015625,0,0.0703125,-0.0078125,0.0390625,-0.0703125,-0.0390625,-0.0234375,0.0234375,0.0078125,-0.0234375,-0.0390625,0.0859375,-0.0078125,0.078125,0.0625,-0.0078125,-0.140625,0.0703125,0,-0.1328125,-0.046875,0.0234375,0.03125,-0.1328125,-0.03125,0.046875,-0.015625,-0.046875,-0.0078125,-0.03125,-0.0234375,-0.015625,-0.0546875,-0.0234375,0.1015625,0.0234375,-0.0078125,0.0078125,0.0234375,0.0078125,-0.015625,-0.0546875,-0.015625,-0.0078125,0.015625,-0.0078125,0.0859375,-0.0546875,0.0078125,-0.0078125,-0.0390625,0,0.046875,0.0390625,-0.0234375,-0.03125,-0.015625,0.0078125,-0.03125,-0.0546875,0,-0.0546875,0.0859375,-0.0546875,-0.0234375,-0.0546875,-0.03125,0.0234375,0.0859375,0.0234375,0.015625,0,-0.0234375,0,-0.0078125,-0.015625,0.015625,0.015625,0,-0.0859375,0.046875,-0.0703125,0.046875,-0.03125,-0.03125,0.0234375,0.078125,-0.0234375,0,-0.0234375,0,0.0390625,-0.015625,-0.0078125,0.0078125,-0.0234375,0.0234375,-0.03125,-0.078125,-0.015625,0.0078125,-0.015625,0.0078125,0.0234375,0.03125,-0.0234375,-0.0078125,0.015625,-0.0078125,0,-0.0078125,-0.015625,0,0.0078125,0.0078125,-0.0625,-0.0234375,-0.03125,-0.015625,-0.046875,0.0078125,0.0078125,-0.015625,0.0234375,-0.0546875,0.0390625,0,0,-0.0390625,-0.03125,-0.0390625,-0.015625,-0.03125,-0.0078125,-0.015625,-0.015625,0.03125,0.015625,0.0390625,-0.015625,-0.046875,-0.0078125,-0.0625,-0.0078125,0.0078125,0,0.0078125,0.03125,-0.0390625,-0.015625,-0.0078125,0,-0.0078125,-0.015625,-0.0703125,0.0234375,-0.03125,-0.0234375,-0.0390625,-0.0234375,-0.03125,-0.0078125,-0.0234375,0.0234375,-0.0234375,-0.0078125,0,0.0078125,-0.0234375,0.0078125,0.0078125,0.0390625,-0.0078125,0,0,-0.015625,-0.0078125,0,-0.0078125,-0.0234375,0,0.078125,0.0078125,-0.0078125,-0.0234375,-0.0078125,-0.0390625,-0.015625,-0.046875,-0.0234375,-0.03125,0.0078125,-0.0390625,-0.015625,-0.015625,0.015625,0.03125,0.0546875,-0.0625,0.0078125,-0.0390625,-0.015625,0.015625,0.0390625,0,-0.0078125,-0.015625,0.0078125,0.015625,0.0234375,0.046875,0,0,0.0078125,-0.0234375,0.0390625,0.0078125,0.015625,-0.0234375,0.0078125,0.0234375,-0.0234375,-0.046875,0.0546875,-0.0390625,0.078125,0,0,-0.0234375,-0.015625,-0.0078125,0.0078125,-0.03125,-0.046875,-0.03125,-0.0390625,-0.03125,-0.03125,-0.03125,0.0078125,0.0078125,0,-0.078125,0.046875,0.0234375,-0.0234375,-0.015625,0.0390625,0.0390625,0.0078125,0.0234375,0,-0.0078125,0.0078125,-0.0546875,0.0078125,0,-0.03125,-0.03125,-0.09375,-0.0078125,-0.03125,-0.0078125,0,-0.0390625,0.0234375,0.03125,0.0546875,0.0234375,0.0078125,0.078125,-0.015625,-0.015625,-0.0078125,-0.03125,-0.0078125,-0.0234375,-0.0078125,0.0625,-0.0390625,-0.0078125,-0.0234375,-0.0390625,0.03125,0.015625,0.0078125,0,0.0859375,0.03125,0,-0.0234375,0.015625,0.03125,-0.0703125,0.0234375,0.015625,-0.03125,0.0078125,0,0.046875,0.078125,-0.0390625,0.0546875,-0.0546875,0.0546875,0.03125,0.0390625,0.015625,-0.0078125,-0.0390625,0.0078125,0.0234375,-0.03125,0.09375,-0.0703125,-0.015625,0,0.09375,0.078125,0.0234375,-0.0390625,0.015625,-0.015625,0.0234375,0.0078125,0.0078125,0,0.0859375,0.0390625,-0.046875,-0.0390625,-0.0625,0.046875,-0.0234375,-0.03125,-0.0703125,-0.0546875,0.0703125,0.0390625,0.03125,0.0234375,0.0546875,0.0234375,-0.0546875,-0.109375,-0.0390625,-0.0234375,-0.015625,-0.0234375,0.0625,0.0390625,-0.0859375,-0.0390625,-0.0234375,0.046875,-0.03125,0.015625,0.0703125,0,-0.0078125,0.03125,0.015625,-0.0234375,-0.0234375,0.015625,0.0078125,0.0078125,0.03125,0.0078125,-0.03125,-0.015625,-0.03125,-0.0078125,-0.0078125,-0.0234375,0.0390625,-0.0078125,0.078125,0,-0.0390625,0.0078125,-0.0078125,-0.0234375,-0.0546875,-0.0078125,0.0078125,-0.0390625,-0.109375,0.0546875,0.0234375,-0.0234375,-0.0234375,-0.0625,0.03125,-0.015625,-0.0078125,0,0,0,0,-0.0078125,0.0078125,0,0.0234375,0.0625,0.0234375,-0.046875,-0.03125,-0.0625,0.03125,-0.0546875,-0.015625,0.03125,-0.0546875,-0.015625,0.0703125,-0.0078125,-0.0546875,-0.046875,-0.0859375,0.0234375,0.1015625,-0.0625,-0.03125,-0.078125,-0.09375,0.0390625,-0.015625,-0.015625,0.1171875,0,0.0078125,0,0,0.0078125,-0.0625,0.0078125,-0.03125,0.015625,0.0390625,0.0703125,0.046875,-0.0078125,0.125,-0.015625,-0.0546875,-0.0078125,-0.015625,0,-0.015625,0.0234375,-0.0390625,-0.0625,0.015625,0.03125,-0.0234375,-0.0078125,-0.03125,-0.0234375,0.0078125,0.0234375,0.0390625,-0.03125,0,-0.015625,-0.03125,-0.015625,0,0.0390625,0.046875,-0.0703125,0,0.0078125,0.0078125,0,-0.0546875,-0.03125,-0.03125,0.0078125,0.0703125,0.0078125,-0.0703125,-0.03125,0.0078125,0.0859375,0.0234375,-0.015625,-0.078125,0.046875,-0.0078125,-0.03125,-0.0078125,0.0234375,0.0234375,0.0234375,0,0,0,0,-0.0078125,0,0,0.0390625,0.015625,-0.046875,-0.03125,0.0390625,-0.015625,0,-0.0234375,-0.0234375,-0.1015625,-0.078125,0.0390625,0,-0.09375,0.015625,0.0078125,0,-0.0078125,-0.015625,0.046875,0.0078125,-0.0390625,-0.046875,0.0078125,-0.0078125,-0.0546875,0.0546875,0.078125,0.0234375,0.015625,-0.0390625,-0.0390625,-0.0703125,-0.03125,-0.0234375,-0.0546875,-0.0390625,0.0546875,-0.046875,-0.046875,0.015625,-0.0078125,-0.03125,-0.078125,-0.0390625,-0.0078125,0.109375,-0.0390625,0,-0.1328125,0.0078125,-0.015625,0.0390625,-0.0078125,-0.03125,-0.078125,-0.0390625,0.1171875,-0.0859375,0.0234375,0.03125,-0.015625,0.015625,-0.0078125,-0.015625,0.0078125,0,0.046875,0.0078125,-0.046875,-0.0390625,-0.0078125,-0.046875,0.0390625,0.015625,0.0078125,-0.046875,-0.0078125,-0.046875,-0.09375,0.0234375,-0.0234375,-0.046875,-0.0234375,0.0546875,0.0078125,-0.046875,0.0234375,-0.0390625,0.0078125,-0.078125,-0.03125,0.0234375,-0.0703125,0.046875,0.0703125,-0.0625,0.1015625,-0.0078125,-0.0625,-0.03125,0.0234375,0.046875,-0.015625,-0.046875,0.015625,-0.0078125,-0.015625,-0.0546875,0,0.0625,0.1015625,0.15625,-0.046875,-0.0078125,-0.03125,-0.0234375,0.109375,0.015625,0.0625,0.109375,-0.0078125,-0.015625,0.015625,0.015625,-0.0078125,-0.0078125,0.1015625,-0.0546875,-0.03125,0.015625,0.0625,0,-0.0703125,-0.0234375,-0.0390625,-0.0859375,0.0078125,-0.0625,-0.0234375,0,-0.046875,-0.03125,-0.046875,-0.0078125,0,-0.0078125,-0.0078125,-0.015625,0.0078125,0.0078125,0.0078125,0.0078125,0.046875,0.0859375,0.0390625,-0.0078125,0.09375,-0.1328125,-0.0625,0.015625,-0.0625,0,-0.0234375,0.015625,-0.0234375,0.0234375,-0.015625,-0.015625,-0.0234375,-0.109375,-0.0234375,0.0390625,-0.0078125,0.0078125,-0.0703125,0.1171875,0.0078125,-0.0625,-0.046875,-0.0078125,0,-0.015625,0.015625,-0.015625,0.015625,-0.015625,-0.015625,0.0078125,-0.015625,-0.0234375,-0.0625,-0.046875,0.0546875,0.03125,-0.0234375,-0.046875,-0.0625,0.09375,-0.0703125,0.03125,-0.0390625,-0.1171875,-0.0546875,-0.046875,0.0078125,-0.03125,0.0078125,0.140625,-0.0078125,-0.15625,0.0703125,-0.1640625,0.046875,-0.0234375,-0.015625,-0.0078125,0.0390625,-0.0234375,0,0.0546875,-0.0703125,-0.0234375,0,-0.0546875,0,0.0625,-0.03125,0.0234375,-0.0234375,-0.0078125,-0.0234375,0,0.046875,0,-0.0234375,0.0078125,-0.0234375,0.0078125,0.03125,0.0078125,0.046875,-0.015625,0.0859375,0.0390625,0.015625,0,0.0390625,-0.015625,-0.0234375,-0.0234375,0.03125,0,0.0625,0.015625,0.015625,0.0078125,0.015625,-0.03125,0.015625,-0.0390625,-0.046875,-0.0703125,0.078125,-0.03125,-0.0390625,-0.03125,-0.0078125,-0.1015625,0.046875,-0.046875,0.0390625,-0.0625,-0.0390625,-0.0078125,0.046875,-0.03125,-0.0703125,0.0546875,-0.0078125,-0.0078125,-0.0078125,-0.0078125,-0.015625,-0.0234375,0.0078125,-0.015625,-0.0078125,-0.0078125,-0.1328125,0.0078125,-0.0078125,0.0078125,-0.0078125,-0.0234375,0.0078125,-0.0390625,0.0703125,-0.0703125,0.0703125,-0.015625,-0.0078125,-0.046875,0,0.078125,-0.046875,0.0234375,-0.0390625,0,-0.03125,-0.0546875,-0.03125,0.03125,-0.0625,0.0390625,0.046875,-0.03125,0.03125,0.03125,0.015625,-0.03125,-0.03125,-0.0859375,-0.0625,-0.0078125,-0.09375,0.0390625,-0.078125,-0.046875,0.046875,-0.0859375,0.0078125,0.1640625,0.015625,-0.0078125,-0.0625,-0.046875,0.09375,-0.0078125,-0.0390625,-0.0234375,-0.0625,-0.0390625,-0.1015625,-0.0234375,0.1640625,0.09375,0.015625,-0.1171875,0.1484375,-0.0859375,0.015625,-0.03125,0.046875,0.0390625,0.0546875,0.015625,-0.0859375,-0.0078125,0.0078125,-0.0078125,-0.015625,-0.03125,-0.03125,-0.0078125,-0.0078125,-0.125,-0.0234375,-0.03125,0.0390625,0.09375,0.0625,0.015625,-0.0625,-0.03125,0.03125,0.03125,0.125,-0.015625,0.0234375,0.0078125,0.0546875,0.0390625,-0.03125,-0.0703125,0.03125,0.0234375,-0.0390625,-0.0625,-0.015625,0.0390625,0,0.0234375,-0.0546875,0.015625,0.03125,0.0078125,0.015625,0.0234375,0.015625,0.03125,0.0234375,-0.0625,0.0546875,-0.03125,0,-0.03125,-0.015625,-0.0546875,0.015625,-0.0234375,-0.03125,-0.015625,-0.0390625,0.0234375,-0.1328125,0,-0.015625,-0.0703125,-0.046875,-0.015625,0.15625,0,0.0234375,0.0390625,0.0078125,0.0078125,-0.0390625,-0.0234375,0.078125,0.03125,-0.0234375,0.0234375,0,-0.0078125,0.0078125,-0.0078125,0.0078125,-0.0078125,0,0.0234375,-0.015625,0.0234375,0.0234375,-0.03125,-0.0390625,-0.0390625,0.0546875,-0.046875,-0.0234375,-0.0078125,-0.0546875,-0.0078125,-0.046875,0.0234375,-0.0078125,0.0234375,0.0390625,-0.0859375,-0.0625,-0.0078125,-0.0390625,-0.03125,0.1328125,-0.015625,-0.0390625,-0.046875,0.03125,0,0.0078125,-0.015625,-0.0078125,0.0078125,-0.0078125,0,0,-0.0078125,0.0234375,-0.046875,0.03125,0.09375,-0.078125,-0.0625,-0.046875,-0.0078125,-0.015625,-0.0234375,-0.078125,-0.078125,-0.0234375,0.03125,0.03125,0.03125,0.0078125,-0.015625,-0.0390625,-0.03125,-0.0859375,-0.078125,0.0546875,0.0390625,-0.0546875,0.0625,-0.046875,0.0078125,-0.015625,-0.0078125,-0.0546875,-0.0625,-0.015625,0.0546875,-0.046875,-0.0078125,0.015625,-0.0078125,-0.0078125,-0.015625,0,-0.0625,0.0234375,-0.0390625,-0.0234375,0.0234375,-0.0390625,-0.0078125,0.03125,-0.015625,0,-0.0703125,-0.046875,0.0078125,-0.0390625,0.0078125,0.0078125,0.0078125,-0.03125,-0.0234375,-0.015625,0.03125,-0.015625,-0.0234375,-0.0234375,0.0546875,0.0390625,-0.015625,0.046875,-0.0234375,-0.03125,-0.015625,-0.0546875,-0.046875,-0.0234375,0.015625,-0.03125,0.0234375,-0.0078125,0,0.0390625,0.0234375,-0.0625,-0.046875,-0.0234375,-0.046875,-0.03125,0.0625,0.0078125,0.1015625,0.0078125,0,0.0078125,-0.015625,-0.0078125,0.0078125,-0.0078125,-0.015625,-0.0078125,0.140625,0.109375,-0.015625,-0.0859375,-0.0703125,-0.0703125,-0.0390625,0.0078125,0.0078125,-0.03125,-0.015625,-0.046875,0.0234375,-0.03125,0.0859375,0.03125,-0.0078125,0.0078125,-0.0546875,-0.0859375,-0.03125,0.0078125,0.046875,0.015625,0.0234375,-0.015625,-0.0234375,0.03125,0.0234375,-0.0546875,-0.0390625,-0.0546875,0.0390625,-0.0234375,-0.0625,0.0234375,-0.0390625,0.0078125,-0.046875,0.0234375,0,0.0390625,0.046875,0.0234375,0,0.0546875,0.0390625,-0.0234375,-0.0078125,-0.0234375,0.03125,-0.0078125,-0.0078125,-0.03125,-0.03125,0.015625,-0.0234375,-0.0703125,-0.09375,0.1015625,-0.015625,-0.0625,0.046875,0.0390625,0,-0.0234375,0.046875,-0.0546875,-0.0234375,-0.0625,-0.0390625,-0.0234375,0.015625,0.0625,0.0625,0.078125,0.046875,0.0703125,-0.03125,-0.09375,0.0234375,-0.0859375,0.0078125,-0.0234375,0.078125,0.0859375,0,0.0390625,0.0703125,0.0078125,0.015625,0.0859375,0.0390625,0.1171875,-0.0703125,-0.0390625,-0.03125,-0.078125,0,0.015625,-0.0625,0.0234375,0.0234375,0,0.0625,0.0625,-0.0078125,-0.0078125,0.046875,-0.046875,0.03125,0.015625,0,0,0.03125,0.015625,0.03125,0.078125,-0.078125,0.015625,0.015625,-0.015625,0.0078125,-0.0390625,0.0234375,-0.03125,0.0390625,-0.03125,-0.015625,-0.0390625,-0.09375,0,0.0234375,0.015625,0.015625,0.0390625,-0.0546875,-0.015625,0,-0.0078125,-0.0234375,0,-0.0390625,0.0390625,0.0078125,-0.0078125,0.0078125,-0.0078125,-0.015625,0.015625,-0.015625,0.015625,0,0.015625,0.046875,-0.0078125,0.03125,-0.078125,-0.078125,-0.0390625,0.015625,0.125,0.03125,0.0234375,0.0234375,-0.0078125,-0.0234375,0,-0.0625,0.015625,0.0078125,-0.03125,-0.0078125,-0.0390625,0.015625,-0.0234375,-0.046875,0.0390625,0,0.0234375,0,0.0078125,-0.0078125,-0.0078125,-0.0078125,0,-0.0078125,-0.0078125,0.0078125,-0.0078125,-0.046875,-0.0234375,-0.0390625,-0.0234375,-0.015625,-0.0546875,0.109375,-0.0625,0,0.0234375,-0.015625,-0.0078125,-0.015625,0.03125,-0.0078125,0.046875,0.09375,0.0390625,-0.03125,-0.03125,0,-0.0234375,-0.0390625,-0.015625,-0.0625,0.0546875,0.015625,-0.03125,-0.0078125,0,-0.015625,-0.015625,-0.0234375,0.0078125,0.0390625,0.0625,-0.0390625,-0.0546875,0.0078125,0.0546875,-0.0078125,0.0546875,0.015625,-0.0625,-0.015625,-0.015625,0,-0.046875,-0.03125,0.0625,0.015625,0.0390625,0.0546875,0.0078125,0,0.0078125,-0.0234375,-0.0078125,0.015625,-0.0078125,-0.0078125,0.015625,0,0,-0.015625,-0.046875,-0.0390625,0,0.03125,-0.0390625,-0.0390625,-0.0234375,0,0,-0.0078125,0.0078125,-0.0703125,-0.0078125,0.0546875,-0.0078125,-0.015625,0,-0.0390625,0.03125,0.03125,0.0078125,0.0234375,-0.03125,-0.09375,-0.0078125,0.0078125,0,0.0078125,-0.0078125,-0.0234375,-0.0078125,-0.0234375,-0.0078125,0.03125,0,0.0078125,-0.015625,0.015625,-0.0234375,-0.03125,0.0390625,0.03125,-0.015625,-0.0234375,0.0234375,-0.03125,-0.0078125,0.0078125,-0.0078125,0.03125,0.03125,-0.0390625,0.0234375,0.015625,0,-0.0703125,-0.0234375,-0.0078125,-0.0078125,0.0859375,-0.0234375,0.0078125,-0.0078125,-0.0625,-0.046875,0.0390625,0,0.0234375,-0.046875,-0.0078125,0.0078125,0.0234375,0,-0.0390625,0.0234375,0.03125,-0.0234375,0.015625,-0.015625,0.03125,-0.03125,0.015625,-0.0703125,-0.0390625,0.0390625,-0.0234375,0.0390625,-0.0546875,0.0234375,0.0546875,-0.015625,-0.015625,0,0.0078125,-0.0234375,-0.046875,-0.0546875,0.0078125,0.03125,-0.0546875,0.0078125,0.015625,0.0234375,-0.0234375,0.0859375,-0.015625,0.046875,0.0390625,-0.0078125,-0.078125,-0.1015625,0.1171875,-0.0390625,-0.0234375,0.0078125,-0.0234375,-0.03125,0,0.0078125,0.03125,0.015625,-0.03125,0.0390625,0.0390625,-0.03125,-0.0546875,0.046875,-0.0234375,-0.0234375,-0.03125,-0.0546875,-0.09375,0.0390625,-0.0234375,-0.0078125,-0.0625,0.015625,-0.0078125,-0.0234375,-0.046875,0.015625,-0.015625,0.046875,-0.0078125,0,-0.0078125,0.015625,0.015625,0.0078125,-0.046875,-0.0078125,0.0234375,-0.0234375,-0.0390625,-0.0234375,0.015625,0.03125,0.0390625,0.03125,-0.015625,0.0078125,0.0078125,-0.03125,0.03125,0,-0.046875,-0.0390625,0.0234375,0,0.0390625,0.0078125,0,0.015625,-0.0625,-0.0234375,0.078125,-0.0078125,-0.0078125,0,0.015625,-0.015625,-0.015625,0.015625,-0.0078125,0,0.0078125,0.015625,-0.0234375,-0.0234375,-0.046875,-0.015625,-0.03125,0,0.015625,0.03125,0,0.0234375,0,-0.03125,-0.0859375,0.0078125,-0.0078125,0,0.015625,0.03125,-0.0078125,0.03125,-0.03125,-0.078125,-0.0625,0.0390625,0.015625,0.015625,0.0078125,0.015625,0,-0.0078125,-0.0078125,-0.0078125,0.0078125,-0.0078125,0,0.03125,-0.046875,0.078125,-0.0546875,-0.078125,0,-0.046875,-0.1015625,0.0078125,-0.015625,-0.0625,-0.015625,0.0078125,0.03125,-0.046875,0.078125,0.09375,-0.046875,-0.015625,0.046875,0.2421875,-0.0390625,-0.0546875,-0.046875,-0.0390625,-0.0859375,-0.0234375,-0.0390625,-0.0546875,-0.0390625,-0.0234375,-0.0234375,-0.03125,-0.0234375,0.0234375,0,-0.0390625,0.0078125,-0.0078125,0,-0.0625,-0.0078125,0.0390625,-0.0078125,0.0234375,-0.0234375,-0.015625,0.0234375,0.0390625,0.09375,0.0703125,-0.0234375,-0.0078125,-0.0546875,0,0.0546875,0,0,0.046875,0.03125,-0.0078125,-0.0078125,-0.0078125,0.0390625,-0.0078125,-0.0078125,-0.0625,-0.046875,0.015625,0,-0.0078125,-0.015625,-0.0390625,0.0703125,0.0234375,-0.0390625,-0.0625,0.0234375,0.0390625,0.0390625,0.015625,-0.015625,-0.015625,0.078125,0.015625,-0.0625,-0.0703125,0.03125,0.03125,0.046875,0,-0.0234375,-0.0078125,0.015625,0.0078125,0,0.0078125,0.0390625,0,0.0078125,-0.0078125,-0.0078125,-0.046875,0.046875,0,0,-0.0234375,-0.0078125,0.015625,-0.015625,-0.0078125,-0.0078125,0.109375,0.0390625,-0.046875,-0.0625,-0.046875,0.03125,-0.03125,0.015625,-0.015625,-0.0078125,0.0703125,-0.03125,-0.0078125,0.0078125,0,-0.0390625,-0.03125,0.0078125,0.015625,-0.0078125,0.0390625,0.015625,0.046875,0.0234375,-0.0234375,-0.0234375,0.0625,-0.015625,-0.03125,0,-0.0078125,0.015625,-0.0234375,0.0234375,0,-0.0390625,-0.0234375,0.1171875,-0.0078125,-0.03125,0.078125,0.0390625,-0.109375,0.1484375,-0.046875,-0.0546875,0.0234375,-0.1015625,-0.0390625,-0.0234375,0,-0.0234375,0,0,-0.0546875,0.078125,-0.0078125,-0.0625,0.0078125,-0.015625,0,0.015625,0.0078125,-0.046875,0.109375,-0.0078125,0,-0.0546875,-0.0390625,-0.0234375,-0.03125,0.046875,0.0703125,0.015625,-0.03125,0.015625,-0.0625,-0.09375,-0.0234375,-0.03125,0,-0.109375,0.078125,0.0859375,-0.0390625,0.0234375,-0.0078125,0.0546875,0.015625,-0.0234375,-0.125,-0.0234375,0.03125,-0.0078125,-0.0703125,-0.0078125,0.0703125,0,0.0078125,-0.1015625,0.0234375,-0.0234375,-0.03125,0.0234375,0.0390625,-0.0390625,0.046875,-0.0546875,0.0390625,0.03125,-0.046875,0.0078125,-0.0078125,0.0390625,0.0078125,0.015625,0.078125,-0.046875,0.015625,-0.0078125,-0.03125,0.0078125,-0.015625,0.0390625,0,-0.0390625,0.1171875,0,-0.046875,0.0390625,0.0234375,0.0078125,0,0.0078125,0.0078125,0.015625,0,0.015625,0.0078125,0,0.0390625,0.046875,-0.046875,0.046875,-0.0234375,-0.0703125,-0.03125,-0.0703125,0.03125,0.0078125,-0.0078125,0.0390625,-0.0390625,-0.046875,-0.0234375,-0.0390625,-0.0234375,-0.0390625,0.0234375,-0.015625,-0.0234375,-0.0078125,-0.03125,-0.03125,0.046875,0.0078125,-0.0234375,-0.0078125,0.0078125,0.0078125,-0.0078125,0,0,0.0078125,-0.015625,-0.0078125,-0.0390625,0.046875,-0.046875,-0.015625,0.0703125,-0.015625,-0.0234375,-0.03125,0.0625,0.0859375,-0.0390625,0.015625,-0.0625,-0.0234375,-0.0078125,-0.0078125,0.0859375,0.0546875,-0.015625,-0.0703125,0.0078125,-0.078125,-0.0546875,-0.0703125,0.109375,0.0625,-0.0390625,-0.015625,0,-0.0234375,0.015625,-0.03125,0,-0.03125,-0.015625,0.0234375,0.0234375,-0.0234375,-0.046875,-0.015625,0.0625,-0.0625,0.0078125,0.0390625,-0.0078125,-0.03125,-0.0234375,-0.0234375,0.0234375,-0.0234375,0,0.0234375,-0.015625,0,0,-0.015625,0.0078125,0.03125,-0.0234375,0.015625,-0.0078125,0.03125,0.03125,0,-0.0390625,0,-0.03125,-0.0546875,0.0390625,0.0234375,-0.0078125,-0.03125,0.0234375,-0.0625,0.0234375,0.03125,0.0703125,-0.03125,-0.0234375,0.046875,-0.0078125,0.0234375,0,0,0.0625,0.0390625,0.0390625,-0.015625,-0.078125,0.015625,-0.0078125,-0.015625,-0.0078125,-0.0078125,0.015625,0.0078125,0,0.0390625,0.0078125,-0.0078125,-0.015625,-0.0078125,-0.015625,-0.0234375,-0.0078125,0,-0.03125,0.0078125,-0.03125,-0.0234375,0.0078125,0.0390625,-0.0234375,-0.03125,0.0234375,0.015625,-0.0546875,-0.015625,0,-0.0390625,-0.0390625,-0.0625,-0.015625,-0.0078125,0.03125,0.03125,-0.015625,-0.0859375,0.015625,-0.046875,0.03125,0.0625,0.0078125,0.1328125,-0.0390625,0.015625,0.015625,-0.0078125,0.0625,-0.0234375,0.0078125,-0.0625,0.0390625,0.015625,0.0078125,0.0546875,-0.0078125,0.0546875,-0.109375,-0.0234375,-0.0234375,-0.0234375,-0.0078125,-0.0390625,-0.0234375,-0.0390625,-0.03125,0.0234375,0.0546875,0,-0.0625,-0.0390625,-0.0078125,-0.015625,-0.0078125,0.0234375,-0.015625,-0.0546875,0.03125,0.0234375,-0.0703125,0.078125,-0.0234375,-0.0234375,-0.03125,-0.0625,0,0.03125,-0.015625,-0.0546875,-0.0234375,-0.015625,-0.0078125,0.015625,-0.046875,0.0078125,0,-0.015625,0.0546875,-0.015625,-0.0234375,-0.0390625,0.0390625,0.0234375,0.03125,-0.03125,0.0078125,-0.09375,0.03125,-0.0546875,0.0078125,-0.0078125,-0.1015625,0.0390625,-0.09375,0.09375,0.0078125,0.0546875,0.0078125,0.0078125,-0.0078125,-0.03125,0.0234375,-0.0078125,-0.0625,0.0234375,-0.0078125,0.0390625,0.015625,0.046875,0,0,0,-0.0234375,0.0390625,-0.0546875,0.03125,-0.015625,-0.046875,0.0234375,0.0703125,-0.0234375,0.0078125,-0.0625,-0.015625,0.0703125,0.0078125,-0.0546875,0.03125,-0.015625,-0.015625,-0.0234375,0,-0.015625,-0.015625,0,-0.0078125,0.0078125,0,-0.0078125,0.0078125,0,0.03125,-0.0546875,0.015625,0.1015625,0.015625,-0.03125,0.0234375,-0.078125,0.0078125,-0.046875,-0.0625,0.0546875,0.03125,0.0546875,-0.015625,0.046875,0.0625,0.015625,0.0078125,0.015625,0.015625,-0.0546875,0.046875,-0.0234375,0.03125,0,-0.0078125,0,0,-0.015625,-0.0078125,-0.0078125,0,0.0078125,0.0078125,-0.0078125,-0.0390625,0.0859375,0,-0.0546875,0,0.0234375,0.0078125,-0.046875,-0.0390625,-0.046875,-0.0859375,0.0078125,-0.046875,-0.0390625,-0.0234375,-0.0546875,0,0.015625,0.0078125,-0.0078125,-0.046875,0.03125,0.015625,-0.0625,-0.03125,0.046875,0.03125,0.0078125,0.015625,0.0234375,-0.0078125,0.015625,0.046875,-0.015625,-0.015625,-0.03125,0.0390625,0.0390625,0.03125,-0.03125,-0.0625,0,0,-0.0625,0,-0.0390625,-0.0703125,0.03125,0,-0.015625,0.0078125,0.0078125,-0.0234375,-0.0078125,-0.0234375,0.0078125,0,-0.015625,0,0.0078125,-0.015625,0.03125,-0.0078125,0.0078125,0.03125,0.03125,-0.0078125,-0.0078125,0.0390625,-0.0078125,-0.015625,0.0078125,0,0.0625,-0.0078125,-0.0546875,-0.0390625,-0.015625,0.0703125,0.0078125,0.0078125,-0.0625,0.0859375,-0.0703125,-0.03125,0.03125,0.0234375,0.0625,-0.0546875,-0.015625,-0.0234375,0,0,0.0078125,0,0.03125,-0.015625,-0.015625,0,0.0078125,-0.0546875,0.0078125,0.0703125,-0.015625,-0.015625,-0.0390625,0.015625,0,0,0.015625,-0.0078125,-0.046875,-0.0234375,-0.0078125,-0.0078125,0.0234375,-0.03125,0.1484375,0.015625,-0.0546875,-0.078125,0.0078125,-0.0546875,-0.046875,-0.03125,0,-0.0078125,-0.0234375,-0.046875,-0.0234375,0.09375,0.015625,0.0078125,0.0078125,-0.0234375,0.03125,-0.078125,-0.0546875,0.0546875,0.078125,0,-0.078125,-0.015625,-0.046875,-0.0234375,-0.015625,-0.0078125,-0.03125,-0.0390625,-0.0546875,0.015625,-0.0390625,0.0234375,-0.046875,-0.0390625,-0.03125,0.015625,0.0625,0.0390625,-0.0390625,-0.015625,0.0234375,0.015625,0.0390625,-0.0390625,0,0.0234375,0.0234375,0,-0.015625,0.015625,-0.046875,0,0.0390625,0.046875,0.015625,-0.0078125,-0.0625,0.0234375,0.0625,-0.015625,0.0390625,-0.03125,0.015625,0,0.03125,-0.0703125,-0.046875,0.0078125,0.015625,0.109375,0.03125,0.015625,-0.0390625,-0.0234375,0.046875,-0.0234375,-0.0390625,0.0234375,0.1171875,0.0078125,-0.046875,-0.03125,-0.0625,0.03125,0.0078125,-0.0234375,-0.0234375,-0.0078125,0.0546875,0.0234375,-0.1015625,0.0234375,-0.0234375,0.0078125,-0.0078125,-0.0625,-0.0234375,-0.0546875,0.0078125,-0.015625,-0.03125,0.0546875,0,0,-0.0078125,-0.0703125,0,0.03125,0,-0.0234375,-0.0234375,0,0,-0.015625,-0.046875,0.015625,-0.015625,0.03125,-0.0234375,-0.03125,-0.0078125,0.046875,0,0.0078125,-0.0078125,0,0.0234375,0.0078125,0,0.0234375,-0.015625,-0.0234375,-0.0078125,-0.0546875,-0.0078125,-0.0078125,-0.0234375,-0.0234375,-0.0390625,0.015625,-0.0078125,0.0546875,0,-0.0078125,0.046875,-0.0390625,-0.015625,0.03125,0.03125,-0.0078125,0.0234375,0.0234375,-0.0078125,-0.015625,-0.0859375,-0.0390625,-0.0625,0.0234375,0.0078125,-0.0078125,0.0078125,0,0.0078125,0.0078125,-0.0078125,0.0078125,0,-0.0078125,-0.015625,-0.0078125,-0.0234375,-0.015625,0.0390625,-0.046875,0.0546875,0,-0.0078125,0.0078125,-0.015625,-0.015625,0.015625,-0.1015625,-0.015625,0.0859375,0.0234375,0.0078125,0,0.03125,-0.0078125,0,-0.0390625,-0.015625,-0.0078125,0.0703125,-0.0078125,-0.015625,0.0234375,0.0078125,0.0078125,0.0546875,0.015625,-0.046875,-0.0078125,-0.015625,0.015625,0.03125,-0.015625,-0.0078125,0.0078125,-0.015625,0.09375,0.0703125,-0.015625,-0.0234375,-0.0234375,-0.015625,0.0078125,0.03125,-0.0078125,0.0390625,0.0234375,0.0078125,-0.015625,0.0078125,-0.015625,-0.015625,-0.03125,-0.015625,0.015625,-0.0078125,-0.0078125,0,-0.0234375,-0.0234375,-0.0078125,-0.03125,0,0,0.0390625,-0.0078125,0.015625,0.0234375,-0.015625,0,-0.046875,-0.015625,0.03125,-0.0234375,-0.015625,-0.046875,0.0625,-0.03125,-0.046875,-0.015625,-0.015625,-0.0703125,-0.0546875,0.0078125,-0.0078125,0,0.0078125,0.0078125,0,-0.015625,-0.0078125,-0.015625,0,0.015625,-0.0234375,-0.015625,0.0078125,0.0390625,0.0078125,0.03125,0.0546875,-0.015625,0.0546875,0.0078125,-0.015625,0.0234375,0.03125,-0.0078125,0.0703125,-0.0234375,-0.015625,-0.0078125,0,0,-0.0078125,-0.109375,0,0.0078125,0.046875,-0.015625,0.0234375,0.0078125,-0.0234375,-0.0234375,-0.046875,-0.0078125,0.0078125,-0.015625,-0.015625,-0.0546875,0.03125,-0.0078125,-0.078125,-0.0390625,-0.015625,-0.046875,-0.0390625,-0.0078125,0,0.0078125,-0.03125,-0.0234375,0.0390625,-0.0390625,0.0078125,-0.0078125,-0.0234375,0.0234375,0.0390625,0,0.0546875,-0.03125,-0.0078125,0.0390625,0.03125,-0.0078125,-0.015625,0.0390625,-0.015625,-0.015625,0.0703125,0.015625,0.0625,-0.03125,0.0078125,-0.0078125,0.015625,-0.015625,-0.015625,-0.0234375,-0.0078125,0.015625,-0.046875,-0.0078125,-0.0234375,-0.0078125,-0.0078125,-0.0234375,-0.03125,-0.0234375,-0.0234375,0.0234375,-0.0234375,-0.015625,0.0390625,-0.046875,-0.0078125,-0.015625,-0.015625,-0.015625,-0.015625,0,0.0390625,0.0390625,-0.015625,0.0078125,-0.0390625,-0.015625,-0.0390625,0.0078125,-0.015625,-0.03125,-0.015625,-0.03125,-0.0625,-0.03125,-0.03125,-0.015625,0.015625,-0.0078125,0.0078125,0.046875,-0.015625,-0.0703125,-0.0546875,-0.03125,0.0234375,-0.0546875,-0.03125,0.046875,-0.03125,-0.0234375,0,-0.0234375,-0.0078125,0.046875,-0.0078125,0.0546875,0.046875,0.046875,-0.015625,-0.046875,0.0078125,0.0390625,0.0078125,-0.0390625,-0.0078125,-0.0078125,0,0,0.0078125,0.0078125,-0.0078125,0.015625,0,-0.0625,-0.015625,-0.0234375,0.0703125,-0.0234375,-0.0078125,-0.0234375,-0.03125,0.0234375,0,0,-0.0234375,0.0078125,-0.0546875,0.03125,-0.015625,-0.046875,0.03125,-0.015625,0.03125,-0.046875,0.0078125,-0.015625,-0.015625,-0.0078125,0.03125,-0.0234375,-0.0078125,-0.015625,-0.0078125,0,0.0078125,0,-0.0078125,0,-0.0078125,-0.0625,-0.015625,0,-0.0390625,-0.09375,-0.0078125,0.09375,0.015625,-0.0390625,0.109375,-0.046875,-0.0390625,-0.0078125,-0.0703125,-0.046875,0.015625,0.0078125,-0.046875,0.0078125,0.0703125,-0.0078125,-0.0546875,-0.0546875,-0.046875,0.0390625,0.03125,0.0390625,0.0078125,-0.0390625,-0.0234375,0.0078125,0.015625,-0.03125,0.0625,0.0078125,0.015625,0.0078125,0.046875,0.03125,-0.1171875,-0.0546875,-0.03125,0.0234375,0.0234375,-0.0078125,-0.0234375,-0.046875,-0.0234375,0.0234375,0.0546875,-0.015625,-0.015625,0,-0.0390625,0.0546875,0.015625,-0.0234375,-0.03125,-0.0078125,-0.0078125,-0.0078125,0.015625,0,-0.0078125,-0.0234375,0.0078125,-0.0234375,0.0234375,0.015625,0.0390625,-0.0078125,0.0078125,-0.0234375,-0.0390625,-0.0078125,-0.046875,-0.015625,-0.078125,0.0703125,0.0625,-0.046875,-0.0234375,0.0390625,-0.0625,0,-0.0546875,-0.046875,0.0078125,0.109375,0,-0.0078125,0,0,0.015625,0.0078125,0,-0.015625,0.015625,0,0.0234375,-0.0625,-0.015625,0.0546875,0.015625,-0.0078125,-0.0390625,-0.015625,-0.0078125,0.0078125,-0.0078125,0.015625,-0.015625,-0.046875,0.03125,-0.0078125,-0.03125,0.0234375,0,-0.0390625,-0.0078125,0.140625,0.0703125,0.0078125,0.046875,0.0859375,-0.0703125,-0.09375,0.0234375,0.046875,0.0625,-0.0859375,0.0234375,0.140625,0.03125,0.015625,0.0546875,-0.0078125,-0.015625,-0.0546875,0.0390625,-0.03125,-0.0546875,0.0859375,-0.0390625,0.03125,0.03125,0.046875,-0.0703125,0.046875,-0.0234375,-0.046875,0.015625,0,-0.0390625,-0.015625,-0.0078125,0.125,0.0078125,0.015625,-0.1640625,-0.0078125,0,0.0546875,-0.0078125,0.0234375,-0.015625,0.0390625,-0.015625,0,-0.0390625,0,0.0078125,0.0234375,0.015625,-0.0625,-0.015625,0.0078125,-0.046875,-0.0546875,-0.0234375,0.0390625,-0.0625,-0.0234375,0,-0.03125,-0.0234375,0.1015625,0.03125,0,-0.0546875,-0.09375,-0.015625,0.0078125,-0.0234375,-0.03125,0.0546875,-0.015625,-0.03125,-0.0625,-0.0390625,0.015625,0.0625,-0.0390625,0.0078125,-0.078125,-0.0234375,-0.0390625,-0.0546875,-0.046875,-0.03125,0.0078125,-0.0234375,-0.0546875,-0.046875,0.015625,-0.015625,-0.015625,0.03125,0.015625,0.0546875,0.0390625,-0.03125,0.015625,0.0078125,-0.03125,0.0390625,-0.046875,0.0078125,0.0078125,0,-0.0078125,-0.015625,0.0234375,-0.0078125,-0.03125,-0.0078125,-0.0390625,0.0078125,0.0625,0.0234375,-0.0078125,-0.03125,-0.0390625,0.015625,0.0078125,0,0.0078125,-0.015625,0.0078125,-0.015625,-0.0078125,0.0078125,-0.0390625,-0.015625,0.0546875,0.015625,0.015625,0,0,0.0078125,0.015625,0.0078125,0.0078125,0.0234375,0.015625,0.0078125,-0.046875,0,0.0234375,0,-0.0078125,-0.015625,0.0703125,0,-0.046875,-0.015625,0,-0.03125,0.0078125,0.0078125,0,0.015625,0.0078125,-0.0078125,-0.0078125,0,0,-0.0078125,0.0234375,-0.015625,-0.03125,-0.0703125,-0.046875,-0.046875,0,0,-0.0078125,0.03125,0.0234375,0.015625,-0.0234375,-0.0859375,0.0625,-0.015625,-0.015625,-0.0234375,0.0859375,0.078125,0.0546875,-0.0234375,-0.03125,-0.0390625,-0.015625,0.015625,0.0234375,-0.0078125,-0.015625,-0.0078125,-0.015625,-0.03125,-0.015625,-0.015625,-0.015625,-0.015625,-0.03125,0.0546875,-0.0234375,-0.015625,0.0234375,0.0546875,-0.0078125,-0.015625,0,0.0390625,0,0.0234375,-0.0234375,-0.0859375,0.0078125,-0.015625,-0.015625,-0.0078125,0.0078125,0,0.0078125,0.015625,0.0078125,-0.0234375,0.015625,-0.0078125,-0.0078125,-0.0078125,0.015625,0.0390625,-0.0078125,-0.0390625,0.0625,0,0.0078125,0.0234375,-0.015625,0.03125,-0.015625,0.0078125,0.0234375,0.0078125,-0.0078125,-0.015625,0,0.015625,-0.078125,0.078125,-0.046875,-0.0234375,-0.03125,-0.03125,-0.0234375,-0.0234375,-0.015625,-0.0234375,0.015625,-0.0078125,-0.0078125,0.015625,0.0078125,-0.0078125,0,0.015625,0,-0.015625,-0.0078125,-0.0390625,-0.015625,0.015625,-0.03125,-0.015625,-0.03125,-0.0234375,-0.0625,0,0.0078125,0,0.0078125,-0.015625,0.015625,0.0390625,0.0546875,0.0234375,0,-0.0546875,0.03125,-0.015625,-0.0546875,-0.0546875,0,0,-0.046875,-0.0546875,0.0234375,0.046875,0,0,0.0390625,-0.015625,-0.03125,-0.015625,0.0078125,-0.09375,-0.03125,-0.015625,-0.078125,-0.0390625,-0.015625,0.0625,0.046875,0.0234375,0.015625,-0.015625,0,-0.0234375,0,0.0078125,-0.1015625,0.1171875,0.0859375,-0.0390625,-0.0234375,-0.015625,-0.0390625,-0.015625,-0.03125,-0.0390625,-0.0234375,-0.0234375,-0.09375,0.03125,0,-0.015625,-0.0390625,0.046875,0,0.0625,0.0234375,-0.09375,0.0546875,-0.0078125,-0.015625,-0.0078125,-0.0234375,-0.0234375,-0.03125,0.0390625,-0.0234375,0.015625,0.015625,0.015625,0.0078125,-0.0078125,-0.0703125,-0.015625,0,0,-0.0234375,-0.0078125,0.015625,-0.0234375,-0.0234375,-0.1015625,-0.0625,0.0234375,0.0859375,0.0625,-0.015625,-0.03125,-0.0078125,-0.0390625,0.0625,-0.0234375,-0.0703125,0.0390625,-0.0390625,0.0078125,-0.0390625,-0.0234375,0,-0.0859375,0,0.0234375,0.015625,0.0703125,-0.015625,0.0234375,0.0546875,-0.046875,0.046875,-0.03125,-0.03125,0.0078125,-0.0078125,-0.0078125,-0.0078125,-0.015625,-0.0078125,-0.0078125,0,0.0390625,0.09375,0,-0.0390625,-0.015625,-0.0234375,0,-0.015625,-0.0078125,0,-0.0234375,0,-0.0078125,0.0078125,-0.0078125,-0.015625,0.0078125,-0.0390625,-0.0078125,0.046875,0.015625,0.03125,-0.015625,0.0234375,-0.03125,-0.015625,-0.03125,0,-0.015625,-0.0703125,0.046875,0.0078125,0.109375,0.015625,-0.0390625,0.015625,-0.0546875,-0.0625,-0.0703125,0.0234375,-0.0703125,0.046875,0.0078125,0,-0.0078125,0.0078125,-0.0078125,0.0078125,0,-0.0078125,0.0078125,-0.046875,0.0234375,-0.0625,-0.046875,-0.015625,0.03125,-0.046875,0.0078125,0.078125,-0.015625,-0.0390625,0,-0.0390625,-0.0390625,0.03125,0,0.0078125,0,0,-0.0546875,-0.0390625,-0.03125,0.203125,-0.0078125,-0.0859375,0.03125,-0.0625,-0.0234375,-0.0078125,-0.046875,-0.0703125,0.09375,-0.0390625,0,0,0,0.0546875,-0.0390625,-0.0234375,0.0234375,-0.0546875,-0.0078125,-0.015625,-0.0390625,-0.0234375,0.0078125,-0.0234375,-0.03125,0,-0.046875,-0.0078125,-0.0234375,-0.0625,-0.03125,0.015625,0.015625,-0.015625,0.015625,0.0078125,-0.0234375,-0.0078125,0.03125,-0.0234375,-0.0078125,-0.0234375,-0.0078125,-0.015625,-0.0390625,-0.046875,0.015625,-0.125,0.015625,0.0390625,0,0.0078125,-0.0546875,-0.0703125,-0.0234375,0.0390625,0.0703125,0.0078125,0.03125,0.0078125,0.0078125,0.0078125,0.046875,0.015625,-0.0234375,0.015625,0.0234375,-0.0078125,-0.0078125,0,0.015625,0.0078125,-0.0078125,-0.0078125,0.03125,-0.0078125,-0.0234375,0,-0.015625,-0.0546875,0.0625,-0.015625,-0.015625,0.0703125,0,-0.0859375,-0.015625,-0.078125,0.1015625,-0.046875,0.09375,0.0546875,0.046875,0,0.015625,-0.0390625,0.03125,-0.015625,-0.046875,0.015625,-0.0234375,-0.078125,-0.0703125,-0.015625,-0.0078125,-0.0546875,-0.0390625,-0.0390625,0.015625,0.03125,-0.078125,-0.015625,0.015625,-0.0078125,-0.015625,-0.046875,-0.046875,-0.03125,-0.0625,0,-0.0234375,0.015625,0.0078125,0.015625,0.0234375,-0.03125,0.0078125,0.0234375,0.046875,-0.03125,-0.015625,-0.0625,-0.046875,0.0234375,-0.1640625,0.09375,0.078125,-0.1171875,0.0390625,-0.0078125,-0.0078125,-0.0078125,-0.015625,0.0703125,-0.0078125,0.0234375,0.0625,-0.0390625,0.03125,0.03125,0.046875,-0.1171875,-0.09375,-0.03125,0.0546875,0.0078125,0.015625,-0.0078125,-0.0234375,-0.0390625,0.078125,-0.109375,-0.046875,0.0078125,0.0078125,0,-0.015625,-0.0234375,-0.0859375,0,0.015625,-0.0078125,0.09375,-0.015625,0.0390625,0.0390625,0.0078125,0.0234375,-0.046875,-0.1640625,-0.046875,0,-0.015625,0.0234375,-0.015625,-0.0234375,-0.015625,-0.0234375,-0.1484375,-0.03125,0.015625,-0.015625,0.0546875,0.0078125,0.0078125,0.0390625,0.0546875,-0.1328125,0.03125,0,0.1328125,0.015625,-0.015625,-0.0703125,0.0078125,0.046875,-0.0625,0.078125,-0.078125,-0.0390625,0.0078125,-0.0625,0.046875,0.09375,-0.0078125,-0.0234375,-0.0625,0.0078125,0.0078125,-0.0625,0.0078125,0.015625,0,-0.0078125,0.0234375,0.0078125,0,-0.015625,-0.015625,-0.015625,0,-0.046875,0.0078125,0.046875,0.03125,0.03125,0.0078125,-0.0390625,-0.0078125,-0.0078125,0.015625,0.0546875,-0.046875,0.046875,0.015625,-0.0859375,-0.0078125,0.0078125,-0.0390625,-0.046875,-0.0078125,0.1015625,0.0078125,-0.015625,-0.015625,-0.0078125,0.015625,0.0078125,0.03125,-0.0078125,0,-0.0078125,0.0078125,0,-0.0078125,-0.0078125,-0.0625,-0.046875,-0.015625,0.1171875,-0.0546875,-0.0234375,0.0390625,0.03125,-0.03125,-0.0859375,0.15625,-0.046875,-0.03125,0.078125,-0.0390625,-0.1328125,-0.015625,0.015625,-0.0078125,-0.0234375,0.0390625,0.03125,0.015625,0.0078125,0.0078125,0.078125,0.0078125,0.015625,0.0703125,0,-0.0625,-0.03125,0,0.03125,0,0.015625,0,0.0078125,-0.03125,-0.015625,-0.0546875,-0.0078125,0.0078125,0.109375,-0.0234375,0.0625,0.0390625,-0.015625,0.0078125,-0.0234375,0.0234375,-0.015625,-0.0078125,0.015625,-0.0234375,0.015625,0,-0.0234375,-0.015625,-0.0078125,0.015625,-0.015625,0.0078125,-0.0234375,-0.046875,-0.046875,0.1171875,0.015625,-0.03125,-0.0078125,-0.0390625,-0.0078125,-0.0078125,-0.0859375,-0.0625,-0.0234375,0.125,-0.0078125,-0.0078125,-0.0078125,0,-0.0390625,0.09375,-0.0078125,0.0078125,0.03125,0.0078125,0.0234375,-0.046875,0.015625,0,-0.015625,0,-0.0234375,0,0,-0.015625,-0.015625,-0.0234375,-0.0234375,-0.0078125,0.0234375,-0.0234375,-0.03125,0.0234375,0.03125,-0.0078125,-0.0078125,-0.0078125,-0.0703125,-0.0078125,0.0078125,-0.0234375,-0.03125,0.0078125,-0.0390625,0.015625,0.046875,-0.0390625,-0.015625,-0.03125,0.078125,-0.0390625,0.078125,-0.046875,0.0078125,0.0390625,-0.0703125,-0.0390625,0.0546875,0.0546875,-0.03125,-0.0234375,0.03125,-0.0078125,0.03125,0.0234375,-0.015625,0.0234375,-0.078125,-0.0078125,-0.03125,0.0390625,-0.015625,0.0234375,-0.1015625,-0.0078125,-0.1015625,0,0.0078125,0.0234375,-0.0859375,-0.0390625,0.0390625,-0.046875,-0.0234375,-0.0859375,0.0546875,0,0.0390625,-0.0234375,-0.0078125,0.0625,0.0625,0.015625,0.03125,0,0.0078125,0,-0.03125,-0.0078125,0,-0.09375,0.015625,-0.03125,0,0.015625,0.0234375,0.0546875,0,0.03125,0.0703125,-0.03125,0.0078125,-0.046875,-0.0625,-0.0546875,0.0078125,0.0078125,-0.015625,0.046875,0,0.0390625,0.03125,-0.0078125,-0.0390625,-0.0625,-0.0078125,-0.078125,-0.0625,-0.015625,-0.0234375,-0.015625,0,0.0546875,0.109375,-0.0234375,-0.015625,-0.0703125,-0.03125,-0.0234375,0.015625,-0.046875,-0.0078125,-0.0078125,0,0.078125,-0.0234375,-0.03125,0.015625,0.0390625,-0.0234375,-0.046875,-0.078125,-0.0625,0.0078125,0.171875,-0.046875,-0.1171875,-0.015625,0.0078125,-0.0078125,0.03125,-0.0546875,0.109375,0.1015625,0.03125,0.0859375,0.0078125,0.0078125,-0.0078125,-0.03125,0.015625,0.0078125,0,0.015625,-0.0078125,0,0,0.0078125,0,0.0625,0.03125,0.046875,-0.03125,0.0078125,0.0078125,-0.0078125,-0.03125,-0.015625,0.0390625,0.0234375,-0.0625,0.0390625,0.0390625,-0.0625,0.015625,-0.015625,-0.0390625,-0.015625,-0.0234375,-0.0625,0.0234375,-0.046875,0.1015625,0,0.0234375,-0.0234375,-0.015625,-0.0078125,-0.0078125,-0.0078125,0.0078125,0.0078125,0.015625,-0.015625,0,0.109375,0.046875,-0.03125,-0.0078125,-0.046875,-0.015625,0.0078125,-0.046875,0,0.03125,0.015625,0.0703125,-0.0546875,0,-0.0703125,-0.0234375,-0.0078125,-0.0078125,-0.03125,-0.046875,0.078125,-0.0703125,-0.015625,0.0234375,0.015625,-0.0234375,-0.015625,-0.0234375,0.0078125,0.0546875,0,-0.0234375,-0.0390625,-0.0078125,-0.03125,-0.0078125,-0.0390625,-0.0390625,0.1015625,-0.0078125,0.015625,0,0,0.03125,-0.03125,-0.0390625,0.015625,-0.0390625,0,-0.0078125,-0.0234375,0.0078125,0.015625,0.015625,0.0234375,-0.03125,-0.0546875,0.015625,0,-0.0078125,0,0.0078125,-0.0078125,0.0546875,-0.0234375,-0.0390625,0.0234375,0.0078125,0.09375,0,-0.015625,-0.015625,0,-0.0546875,0.0703125,-0.0625,0.0234375,0.0546875,-0.0234375,-0.015625,-0.0625,0.015625,0.0703125,-0.0078125,-0.046875,-0.0546875,-0.0234375,-0.015625,-0.015625,-0.0234375,-0.0078125,0,0.015625,-0.015625,-0.015625,0.015625,0,0.015625,0.015625,0.046875,-0.0625,0,0,0.0078125,-0.0078125,0.015625,-0.0390625,-0.0078125,-0.0234375,0,-0.0859375,0.0625,0.0390625,-0.0546875,-0.0078125,-0.03125,-0.0078125,-0.046875,0.03125,0.0625,-0.078125,-0.046875,0.015625,-0.0234375,-0.0390625,-0.0234375,0.0234375,-0.109375,0.0703125,-0.0078125,0.0078125,0.0546875,-0.0390625,-0.03125,-0.015625,-0.0625,-0.0234375,0.0234375,0.0234375,-0.078125,-0.046875,-0.03125,-0.0546875,0,0.0625,0.078125,0.0078125,-0.078125,0,0.03125,-0.0234375,-0.0390625,0.0078125,0.0390625,-0.046875,-0.0078125,-0.0234375,-0.0390625,-0.0859375,0,-0.0546875,0,-0.0390625,0.0078125,0.015625,-0.046875,0,0.0546875,-0.015625,-0.015625,0,0.0078125,-0.0546875,-0.046875,-0.0703125,0.0390625,0.1171875,-0.015625,-0.015625,-0.015625,0.0234375,0.0234375,-0.015625,0.0390625,-0.046875,-0.0703125,-0.03125,-0.0234375,0.015625,-0.015625,0.109375,-0.0625,0.0859375,-0.0234375,-0.0234375,-0.0078125,-0.0234375,-0.015625,0.0859375,-0.1328125,-0.015625,0.078125,0.0390625,0.0234375,-0.0078125,0.03125,-0.0390625,0.0703125,0.046875,-0.0859375,0.0703125,-0.09375,0.0625,0.0078125,-0.0234375,-0.015625,0.046875,0.0234375,0.0625,0,-0.0703125,0.0078125,-0.0234375,0,-0.015625,0.0078125,0,0.03125,0.0625,-0.0390625,-0.03125,-0.015625,-0.0390625,-0.0078125,-0.03125,0.109375,-0.046875,0.0234375,0.046875,0.0546875,-0.1171875,-0.015625,-0.0078125,-0.0078125,-0.0078125,0,0,0,-0.015625,-0.0078125,-0.0078125,0.015625,0.0546875,0.0390625,0.0234375,-0.046875,-0.109375,-0.0546875,0.0078125,0,-0.0234375,-0.03125,-0.03125,0.046875,-0.0078125,-0.03125,-0.0078125,-0.0234375,0.0390625,0.0703125,0.0234375,0.0078125,-0.0234375,0,-0.1015625,-0.0390625,-0.0078125,0.0234375,-0.078125,0.0078125,0.015625,0.015625,0,-0.0078125,-0.0078125,-0.0078125,-0.0078125,0,-0.0390625,-0.0703125,-0.0390625,0.0234375,-0.0859375,0.0625,-0.03125,0.03125,0.0546875,-0.03125,0,-0.03125,0,0.0234375,0.0078125,0.03125,0.0078125,0.0390625,0.0703125,0.03125,0.0078125,-0.078125,-0.0859375,-0.046875,0.03125,0.03125,-0.0234375,-0.0625,0.0390625,0.03125,-0.0234375,-0.046875,0.0625,-0.0234375,0.0703125,-0.0234375,0.0078125,-0.0078125,-0.0234375,-0.0625,0.0546875,-0.03125,0.015625,-0.109375,0.015625,0,-0.0078125,-0.03125,-0.015625,-0.03125,-0.0546875,-0.03125,0,-0.0078125,0.0234375,-0.0078125,-0.0078125,0.015625,0.0078125,0,-0.03125,0,0.03125,-0.015625,0.046875,0.0078125,-0.0625,-0.03125,-0.0390625,-0.015625,0,-0.046875,-0.0703125,0.03125,-0.0859375,0.015625,-0.0703125,-0.03125,0.046875,0,0.0078125,-0.0078125,0.015625,-0.0546875,0.0625,-0.0546875,0,-0.03125,0.0390625,-0.109375,0,0.0078125,0.0078125,-0.0078125,-0.015625,0.0078125,0.015625,0.03125,0.015625,-0.015625,-0.015625,-0.015625,-0.046875,0,-0.0390625,-0.03125,0.0390625,0.0390625,0.03125,-0.03125,0.0625,0.0078125,-0.0234375,0.0234375,-0.046875,0.0390625,0.0390625,0,0.0234375,-0.0078125,0.0078125,-0.078125,-0.015625,0.0390625,0.015625,-0.03125,-0.0390625,0.09375,0.0078125,-0.125,-0.0078125,-0.1015625,-0.0078125,-0.078125,-0.0234375,-0.03125,-0.0390625,-0.0625,-0.0234375,-0.09375,0.015625,0.0625,0.1015625,0.015625,0.0390625,0.0234375,0,0.0078125,-0.0390625,-0.0859375,0.0078125,-0.0390625,-0.015625,0.03125,-0.0234375,0.078125,-0.0234375,0.03125,-0.0078125,-0.046875,0.015625,-0.0390625,-0.0078125,0.0234375,-0.015625,-0.03125,-0.0078125,-0.0234375,0.015625,0.03125,0.0234375,0,0.0625,0.03125,-0.078125,0.03125,-0.03125,-0.0546875,-0.0078125,0.0234375,-0.0078125,-0.046875,0.0546875,-0.0234375,-0.03125,-0.0390625,0.0234375,0.1171875,-0.0078125,0.15625,0.0078125,0.0234375,-0.0078125,0.078125,-0.03125,-0.078125,-0.0234375,-0.09375,0.015625,0.046875,-0.0390625,0.0625,0.046875,-0.0078125,-0.0078125,-0.09375,0.015625,0.03125,-0.0234375,0.0703125,-0.0546875,-0.015625,-0.0078125,0.078125,-0.0625,0.0703125,-0.0234375,0.0859375,-0.03125,-0.03125,0.046875,-0.0234375,-0.0234375,-0.015625,0.0078125,0.0859375,0.015625,0.046875,-0.015625,-0.0546875,0.015625,-0.0390625,0.015625,-0.0234375,0.125,0.0234375,0.0234375,-0.0234375,-0.1328125,-0.0078125,-0.03125,-0.0078125,-0.015625,0.0078125,0.03125,0,0,-0.015625,-0.0078125,0.0078125,0.0078125,-0.0078125,0,-0.0546875,-0.0078125,-0.03125,0.015625,-0.046875,0.03125,0.015625,0.0625,0.0078125,0,0.0234375,0,-0.015625,-0.015625,0.0078125,0.0546875,0.0078125,-0.0234375,0.03125,-0.015625,0.015625,0.046875,0.0859375,-0.0078125,-0.0625,-0.0078125,0.0078125,0,-0.015625,-0.0078125,-0.015625,-0.0078125,-0.0078125,0.0078125,0.0078125,-0.0078125,-0.0546875,0.0078125,0.078125,-0.0390625,-0.078125,0.078125,-0.0234375,0.078125,0.0625,0.0703125,0.078125,-0.0390625,-0.078125,-0.1171875,-0.046875,-0.0390625,-0.0390625,0.0859375,-0.0078125,0.0234375,-0.046875,0.0390625,0.0234375,0,0.015625,-0.015625,-0.0390625,0.0078125,0.015625,-0.0234375,-0.0234375,0.0546875,0.015625,0.046875,0.03125,0.0859375,0.078125,0.078125,0.015625,-0.0234375,0.0390625,-0.03125,-0.046875,-0.0546875,0.015625,0.0234375,0,-0.0234375,-0.0078125,-0.015625,0.0078125,0.03125,0,0.015625,-0.0390625,-0.015625,0,-0.0078125,-0.0234375,-0.015625,-0.0078125,0,-0.03125,0,-0.0078125,0.015625,0,0.0234375,0.0234375,0.0859375,0,0.0859375,0,0.03125,-0.0390625,-0.0625,-0.078125,-0.046875,0,0.03125,-0.0078125,-0.078125,0.0234375,-0.0078125,0.03125,0.0703125,-0.0078125,-0.0390625,0,0.015625,0.015625,-0.0078125,0.0078125,0.0234375,0.015625,-0.0078125,0,-0.0078125,-0.03125,-0.015625,-0.0234375,-0.0078125,0.015625,-0.0234375,0.0234375,-0.0390625,-0.0078125,-0.0625,0.015625,-0.0234375,0.0703125,-0.046875,-0.0234375,0.046875,-0.0078125,0.0625,0.015625,0.015625,-0.03125,-0.015625,0,0.015625,0.046875,-0.0234375,0.0234375,0.03125,0.046875,0.0390625,0.078125,-0.078125,0.0859375,0,0.0390625,0.015625,0.046875,-0.0546875,0.0078125,-0.0078125,-0.1171875,0.0234375,0.0234375,-0.03125,0.03125,0.0625,-0.0234375,0.078125,-0.0078125,-0.0078125,0.0234375,0.0078125,-0.0234375,0.03125,0.015625,-0.015625,-0.0390625,-0.0859375,0.1015625,-0.0546875,0.0625,-0.03125,0.046875,0.015625,0.0078125,-0.015625,-0.046875,-0.0859375,-0.0859375,-0.0546875,-0.0625,-0.015625,0.0234375,0,0.0234375,0.0234375,0.015625,-0.0703125,-0.0390625,-0.09375,-0.0078125,0.0078125,-0.0078125,0,-0.0078125,-0.015625,0.0234375,-0.0390625,-0.03125,-0.1015625,0.046875,-0.0859375,0.03125,-0.0078125,-0.0390625,-0.0234375,-0.0390625,-0.015625,-0.0625,-0.015625,-0.015625,0.0078125,0,-0.0546875,0.0703125,0,0.0078125,0.1328125,0.0234375,0.0234375,0.046875,-0.0390625,0.0078125,0.0390625,-0.015625,-0.0703125,-0.03125,0.0234375,0.046875,0.03125,-0.015625,0,-0.03125,-0.015625,-0.0625,0.0390625,0.078125,0.0078125,-0.0078125,-0.0703125,-0.0546875,-0.046875,-0.046875,-0.03125,-0.0625,0.0078125,-0.0390625,-0.03125,0.03125,-0.0234375,-0.0234375,0.140625,-0.046875,-0.0078125,0,-0.0078125,0,-0.0078125,0,-0.0078125,0.015625,0.0078125,0,-0.0078125,0.0078125,0.0546875,0.0390625,-0.0703125,0.0703125,0,-0.0390625,-0.046875,0.0546875,-0.0625,0.0234375,0.0703125,-0.0078125,0.0625,-0.0546875,-0.03125,-0.0546875,-0.015625,-0.0078125,0.0078125,-0.0625,-0.015625,-0.078125,0.0390625,0.109375,0.046875,-0.0078125,-0.0078125,-0.0078125,-0.0078125,0.0078125,0,0,0.0078125,-0.0078125,0,0.0546875,0.046875,0.0859375,-0.015625,-0.046875,-0.0546875,0.03125,-0.015625,0.03125,0.0078125,-0.078125,-0.046875,-0.03125,-0.09375,0.0390625,0.015625,0.0390625,-0.0078125,-0.0546875,0.03125,0,0.015625,-0.0234375,-0.0078125,0.03125,0.0234375,-0.0234375,0.046875,-0.0234375,0.03125,0.0078125,0.0078125,0.03125,0,0.03125,0.0078125,-0.046875,0.03125,-0.0625,-0.0234375,0.015625,-0.015625,-0.0078125,-0.03125,0.015625,0.0625,-0.015625,-0.0546875,0,-0.0234375,-0.0390625,0.046875,0.0078125,-0.03125,0.046875,-0.015625,-0.03125,-0.03125,0.03125,-0.0078125,-0.0390625,0,0.0078125,0.0390625,0.03125,0.0078125,-0.03125,-0.0234375,-0.0703125,0.015625,0,0.03125,-0.015625,0.0078125,0.03125,0.03125,-0.0078125,0.0234375,-0.0546875,-0.03125,0,-0.1171875,-0.0078125,-0.015625,0,0.0546875,0.03125,0.0625,-0.0390625,0,0,-0.015625,0,0.0078125,0.0078125,0.015625,0,0,0.0234375,0.0625,-0.0546875,0.0078125,-0.015625,0.0234375,-0.03125,-0.0625,0.0234375,-0.046875,0.0078125,-0.0625,-0.03125,0.015625,0.078125,0.0078125,0,0.015625,-0.0078125,-0.0546875,-0.0546875,-0.0234375,0.046875,0,-0.0625,0.0390625,-0.0234375,-0.0703125,0.015625,0.0625,-0.0625,-0.03125,-0.0625,0.015625,0.0234375,0.109375,0.015625,0.0625,-0.03125,0,-0.03125,0.0390625,0.015625,0.015625,0.03125,0.015625,-0.0546875,0.09375,0.015625,0,0.015625,0.0078125,0,-0.015625,-0.0234375,-0.0390625,0,0.03125,-0.03125,0.125,0.015625,0.015625,-0.0859375,0.046875,0.0234375,0.03125,0.0078125,-0.03125,0.0390625,-0.0390625,-0.0234375,0.03125,0.0546875,0.0078125,0.015625,-0.046875,0.0703125,-0.0625,-0.0078125,-0.0078125,-0.0078125,-0.0078125,0.046875,0.046875,0,-0.109375,-0.015625,0.0078125,0.015625,-0.046875,-0.1015625,0.125,-0.015625,-0.015625,-0.078125,0.0234375,0,0.0234375,0.03125,-0.046875,0.0390625,0.046875,0.0078125,0.03125,0,-0.0546875,-0.03125,-0.03125,0.046875,0.0234375,-0.015625,0.046875,-0.03125,0.0546875,-0.0703125,-0.015625,-0.03125,-0.0078125,-0.078125,0.0546875,-0.0859375,-0.0078125,-0.0546875,0.0546875,0.0625,-0.0078125,-0.015625,-0.0078125,-0.0390625,-0.0390625,0.0546875,-0.0234375,-0.015625,0.0703125,0.0078125,0.015625,0.0703125,0,-0.0625,-0.0625,0.0078125,-0.0078125,-0.03125,-0.03125,0.0078125,0.0078125,-0.015625,0.0078125,0.015625,0,-0.0078125,0,0.0078125,-0.0078125,-0.0234375,-0.046875,-0.0390625,0.0234375,-0.0390625,0.015625,0.0390625,-0.0390625,0.03125,0,-0.046875,-0.03125,-0.0625,-0.0625,0.015625,0.0234375,0.0078125,-0.0859375,0.0546875,-0.0234375,0.078125,0.0859375,-0.0625,0.0234375,-0.1015625,-0.0390625,0,0,-0.0078125,0,0,-0.0078125,0.0078125,-0.015625,0,0,-0.078125,-0.078125,0.109375,-0.015625,-0.0625,0.1015625,0.015625,0.0390625,-0.0234375,-0.078125,-0.0703125,0.015625,0.0078125,0.015625,0.046875,0,0.0234375,-0.09375,0,-0.0234375,0,0.0546875,-0.0625,-0.0546875,-0.015625,-0.046875,0.046875,0,0,-0.046875,-0.0078125,-0.015625,-0.0234375,0.0390625,-0.046875,0.03125,-0.0078125,-0.03125,-0.03125,0.046875,0,0.0078125,-0.015625,-0.046875,0.0546875,0.015625,-0.0390625,0.0078125,-0.03125,0.0234375,-0.0234375,-0.015625,0.046875,-0.0078125,-0.015625,0.0234375,0.0703125,0.03125,-0.03125,0.015625,0.015625,0.015625,0,0.03125,-0.0078125,0.0859375,0.0390625,0.015625,-0.0390625,-0.0078125,-0.0234375,0.015625,-0.046875,-0.0078125,-0.0859375,-0.0625,0.0234375,-0.0625,0.0234375,-0.0078125,-0.0078125,-0.046875,-0.0390625,0,0.0703125,-0.0625,0.0390625,-0.046875,-0.0234375,-0.0234375,-0.0234375,0.0078125,0.0234375,-0.0078125,0,0.0078125,-0.0078125,-0.0078125,0.0234375,0.0546875,-0.0234375,-0.0390625,-0.0546875,0.0078125,-0.0078125,0.0390625,0.0234375,-0.0390625,-0.0078125,-0.046875,0.0234375,-0.0390625,0.0625,0.015625,0.0234375,0.03125,-0.0234375,-0.078125,-0.078125,-0.0234375,0.0625,0.0078125,-0.078125,-0.0859375,-0.078125,0.0234375,0.0625,-0.015625,0.0078125,-0.015625,0.0546875,0.0390625,-0.046875,0.015625,-0.0390625,-0.046875,-0.03125,0.0703125,-0.0234375,0.0546875,-0.0703125,-0.0546875,-0.0390625,-0.015625,0.0390625,-0.0078125,0.0078125,-0.046875,-0.046875,0,-0.0078125,0.015625,-0.0390625,0.015625,0.0234375,-0.015625,-0.1171875,0,0.0234375,-0.0625,0.03125,-0.03125,0.03125,-0.0234375,-0.0625,-0.0546875,0.0078125,0.015625,-0.0078125,-0.03125,0.0546875,0.0546875,0.09375,-0.0234375,-0.0546875,-0.046875,-0.046875,-0.0546875,-0.0625,-0.0546875,-0.0234375,-0.03125,0.078125,0.125,0.0078125,0,0,0.0390625,0.046875,0.015625,-0.0078125,0.1015625,0,-0.1015625,-0.0390625,0,-0.0546875,0.0078125,0.0078125,-0.03125,-0.015625,-0.0546875,0.0390625,0.03125,-0.078125,-0.0390625,0.109375,0,0.015625,0.0546875,-0.0625,0.015625,0.0703125,-0.015625,-0.046875,0.015625,0.03125,-0.0078125,-0.0234375,0.015625,0.015625,0.015625,0.015625,-0.03125,0.015625,-0.0234375,0.015625,-0.0078125,-0.140625,0.03125,-0.0234375,-0.046875,0.0234375,-0.03125,-0.03125,-0.09375,0.015625,-0.0390625,-0.015625,-0.0625,0.0546875,0.0625,0,-0.0078125,-0.015625,0.0234375,0.0078125,-0.0078125,-0.015625,0.0078125,0,0.0234375,0.015625,0.046875,0.0078125,-0.1171875,-0.078125,-0.015625,0.0546875,0.046875,0.015625,0.0390625,0.03125,0.0078125,-0.046875,-0.0234375,-0.0234375,-0.015625,0,0.0703125,0.0390625,-0.0703125,-0.046875,-0.0390625,0.09375,0.015625,-0.03125,-0.0390625,-0.0078125,-0.0078125,0.0078125,0.015625,0,-0.0078125,0.0078125,0.0078125,0,-0.0234375,-0.0859375,0.0234375,-0.03125,0.0234375,-0.03125,0.015625,0,0.0703125,-0.0234375,0.1171875,0.015625,-0.0078125,-0.0625,-0.0234375,0.1015625,0.078125,0.1484375,0.03125,-0.0703125,0.0859375,0,-0.1015625,-0.0546875,-0.0703125,0.1015625,0.0390625,0.0078125,0.0390625,0,0.0234375,-0.046875,-0.015625,-0.0703125,0.0078125,0,-0.0703125,-0.0234375,0.078125,-0.0234375,0.03125,0.0546875,-0.03125,0.0078125,0.0234375,0,-0.015625,0.0703125,0.03125,-0.0234375,0.09375,0,-0.015625,0.0078125,0.0390625,-0.0390625,0.078125,-0.0234375,-0.0546875,0.0234375,-0.0078125,0.0390625,0.03125,-0.0234375,-0.0546875,0,-0.0234375,-0.015625,0.015625,0.0078125,-0.046875,-0.046875,-0.0390625,0.0703125,-0.0078125,0.03125,-0.0078125,0.0078125,-0.0234375,-0.0546875,-0.0625,-0.0390625,0.0546875,-0.015625,-0.0234375,0.015625,-0.109375,0.0234375,-0.0390625,-0.0390625,0,-0.0234375,-0.015625,-0.015625,0,0,0.0078125,-0.0234375,-0.0078125,-0.0234375,0.0390625,0.1015625,-0.0234375,-0.015625,0.078125,-0.0390625,-0.078125,0.015625,-0.0546875,-0.015625,-0.03125,-0.0390625,-0.0234375,0.0390625,0.0234375,0.0234375,0,-0.0078125,0.0390625,0.0078125,-0.046875,-0.078125,0.0546875,-0.0390625,-0.03125,0.0859375,-0.0078125,-0.015625,-0.0546875,-0.078125,-0.0703125,-0.046875,-0.0390625,-0.1015625,0.015625,0.0078125,-0.0234375,0.0546875,-0.0390625,0.0078125,0.0234375,-0.0546875,0.0234375,-0.0078125,-0.0078125,-0.0390625,0.0078125,0.0546875,-0.0625,0.0390625,0.1015625,0.0546875,0.0390625,-0.0859375,0.0625,-0.015625,0.0078125,-0.0703125,-0.0859375,0.1015625,-0.1171875,-0.0625,0.0234375,-0.0078125,-0.0390625,0.0234375,0.0390625,0,0.015625,-0.0390625,-0.03125,0.015625,-0.0078125,0,0.0234375,0.0625,0.0859375,0.109375,0.015625,0.0234375,0.03125,-0.0078125,0.0546875,-0.0625,0.0078125,0,-0.03125,-0.0234375,0.0390625,0.0859375,0.0390625,0.0703125,-0.078125,-0.046875,-0.09375,-0.0546875,0.03125,-0.0234375,0,0.0234375,0.0546875,-0.078125,-0.0859375,-0.09375,-0.1015625,0.03125,-0.0078125,0.0625,-0.046875,0.109375,0,-0.09375,0.0625,0.0703125,0.046875,-0.03125,0.078125,0.015625,-0.0234375,-0.0078125,-0.0234375,-0.0390625,0.09375,0.015625,0.03125,0.0390625,0.0546875,-0.015625,-0.015625,0.0078125,-0.0390625,0.046875,-0.0234375,0.03125,0.078125,0.0078125,-0.0390625,-0.046875,0.0078125,0,0.046875,0.015625,-0.015625,-0.0078125,-0.0078125,0.0078125,0,-0.0078125,-0.015625,0,-0.0078125,-0.015625,-0.0625,0.03125,0.015625,-0.1015625,0,0.0078125,0.03125,0.0546875,-0.0078125,-0.015625,-0.125,0.0078125,-0.03125,0.0546875,-0.0234375,-0.015625,0,-0.015625,0.078125,0.015625,-0.0078125,0.0390625,0.0390625,-0.0234375,-0.15625,-0.0625,-0.0078125,0.0078125,0,0,0,-0.0078125,-0.0078125,0,-0.0078125,-0.0078125,0.0703125,-0.0078125,-0.0234375,0.015625,-0.046875,-0.015625,-0.0390625,0.0859375,-0.0390625,-0.0390625,-0.078125,0,-0.015625,0.0078125,-0.03125,0.0625,-0.0078125,-0.0078125,-0.0234375,-0.0703125,-0.0078125,-0.0234375,0.0625,-0.015625,0.0234375,-0.078125,-0.015625,-0.0234375,-0.0078125,0.0078125,-0.0390625,-0.015625,0.0078125,0.0546875,-0.015625,0.0234375,0,0.015625,0.0078125,0.078125,-0.0546875,-0.015625,0.0234375,0.0078125,-0.0390625,-0.0078125,-0.015625,-0.015625,-0.03125,-0.03125,-0.0078125,0.0078125,-0.03125,-0.015625,0.0390625,0.0078125,0,0,0.015625,-0.0078125,0.0078125,0.015625,0,-0.0078125,0.0078125,-0.0078125,-0.0625,0.0234375,0,-0.046875,0.0078125,-0.015625,0.015625,0,-0.03125,-0.0078125,0.0078125,-0.0078125,0.0078125,-0.0234375,-0.0234375,0.1015625,-0.015625,-0.0546875,-0.0234375,-0.0703125,-0.046875,-0.0390625,-0.0390625,-0.015625,-0.015625,-0.0078125,-0.0078125,-0.015625,0.0078125,-0.015625,0.0078125,-0.015625,0,0.0078125,-0.015625,0.015625,-0.015625,-0.0234375,-0.0078125,0,0.0234375,0,-0.0078125,0.0234375,0,-0.0078125,-0.0234375,-0.03125,0,0.015625,-0.0234375,-0.03125,0,0.015625,-0.0625,-0.0546875,-0.0234375,0.0078125,-0.015625,-0.0078125,0.0703125,0.015625,-0.0625,0.0234375,-0.0546875,-0.0546875,-0.015625,-0.0234375,-0.0078125,0.03125,-0.0234375,-0.0078125,0.0234375,-0.046875,-0.0078125,0.0859375,0.015625,0.0078125,-0.015625,0.0625,0.0078125,-0.046875,-0.015625,-0.0078125,-0.015625,0.0234375,-0.0078125,-0.0078125,0.0234375,-0.015625,-0.1171875,0.078125,-0.0234375,-0.109375,0.0078125,0,0.0390625,0.015625,-0.015625,0.015625,-0.0078125,0.0078125,0.015625,0.0390625,0.015625,-0.03125,0.0234375,-0.0078125,0.03125,-0.0078125,-0.0234375,-0.0625,0,0,0.03125,0.015625,-0.015625,0.0390625,0.03125,-0.0390625,-0.03125,-0.0078125,0.0078125,0.015625,-0.0078125,-0.0546875,0.0625,0.03125,0.0078125,-0.0234375,-0.0625,-0.0234375,0.125,0.1015625,-0.0078125,0.046875,-0.0234375,-0.015625,0.015625,0,-0.0078125,-0.0234375,-0.03125,-0.015625,-0.015625,-0.015625,-0.015625,-0.03125,0.0234375,-0.03125,0,0.03125,-0.0078125,-0.0859375,-0.015625,-0.015625,0.0078125,-0.015625,-0.0078125,-0.0078125,0.0234375,-0.0234375,-0.015625,-0.0859375,-0.0546875,-0.0234375,0.0078125,-0.0078125,0.0703125,0.09375,0.078125,-0.0390625,-0.0390625,0.015625,-0.0078125,-0.03125,-0.0078125,0.0078125,-0.0078125,0,-0.0078125,-0.015625,0.0078125,-0.0078125,0.015625,0.015625,0.015625,0.078125,-0.015625,-0.015625,-0.0703125,-0.09375,0,0.0546875,0.109375,-0.0234375,-0.015625,0.0625,-0.0234375,0.03125,-0.0390625,0.0234375,-0.0078125,-0.0234375,0.0078125,0.0234375,-0.0078125,0.078125,-0.0078125,0.078125,-0.015625,-0.03125,-0.015625,0,0,0.0078125,0,-0.0078125,0.0078125,-0.0078125,0.0078125,0.0078125,0.015625,-0.015625,-0.0078125,-0.0078125,-0.0625,-0.09375,-0.0390625,0.0234375,-0.0078125,0.0234375,0.0078125,0.0625,-0.0390625,-0.0234375,0.03125,-0.0390625,-0.015625,0.03125,-0.0234375,0.046875,-0.03125,-0.015625,0.03125,-0.0078125,-0.015625,-0.046875,-0.0703125,0.03125,0.0078125,-0.0078125,-0.0390625,0.015625,-0.0234375,-0.0234375,-0.0234375,0.0234375,0.0234375,-0.046875,-0.0234375,-0.0546875,0.0078125,-0.0390625,-0.0234375,0.015625,-0.0703125,0.0078125,0.0078125,0.0546875,0,-0.015625,0,-0.015625,0.03125,0.0234375,0,0.03125,-0.0078125,-0.0078125,0.0234375,0.015625,-0.0234375,-0.0234375,0.0234375,-0.015625,-0.0234375,-0.0234375,-0.015625,0.0078125,-0.0078125,-0.015625,-0.0625,0.0234375,0.1640625,-0.046875,0.125,-0.046875,-0.0703125,-0.078125,-0.0078125,-0.0625,0.015625,0.0078125,-0.046875,0.03125,-0.015625,-0.015625,0.0390625,-0.03125,0.046875,-0.0625,0.0234375,0.0078125,0.0078125,-0.0078125,0,0,0,0,-0.0234375,-0.0390625,-0.015625,-0.0234375,-0.015625,0.0234375,-0.0390625,-0.015625,0.0390625,0.0078125,0.09375,-0.015625,0.0078125,0.015625,0.0390625,-0.0234375,-0.0390625,-0.046875,0.03125,-0.0078125,0.0078125,-0.0625,-0.0234375,-0.1015625,-0.0625,-0.046875,0.0234375,0.125,0.03125,-0.03125,-0.0625,0.0390625,-0.0078125,0.09375,-0.0234375,-0.046875,0,0.046875,0.015625,-0.0078125,-0.03125,0.03125,-0.03125,-0.0390625,0.046875,0,0.078125,0.03125,0.0625,-0.015625,-0.0703125,-0.0234375,-0.0078125,0.0390625,-0.0234375,-0.0546875,-0.0546875,-0.0234375,-0.0078125,0.0078125,-0.03125,-0.0390625,0,0.15625,-0.0390625,0.015625,-0.0625,-0.0390625,-0.0078125,-0.015625,-0.03125,0.03125,0.1015625,0.0390625,0.03125,-0.0234375,0.0078125,-0.0546875,0,-0.03125,-0.0078125,-0.0390625,0,0.046875,0.03125,-0.0234375,0.0078125,0,-0.0390625,-0.0234375,-0.0390625,0.0078125,-0.1875,0.0078125,-0.0234375,0.0234375,0.0390625,-0.046875,-0.0078125,-0.015625,0.0546875,-0.0546875,0.03125,-0.046875,-0.0234375,-0.015625,0.0234375,-0.0234375,-0.0078125,0.0546875,-0.03125,0.03125,-0.03125,-0.0703125,-0.0859375,-0.015625,0.0078125,-0.046875,0.03125,-0.1015625,-0.0390625,0.0078125,-0.015625,0.0390625,-0.0078125,0.0703125,0.0546875,-0.046875,0.0078125,0.0390625,0.015625,0.0390625,0,-0.0390625,-0.078125,-0.03125,-0.015625,-0.015625,0.03125,-0.046875,-0.0390625,0.0078125,-0.0703125,-0.0390625,-0.0546875,0.0078125,0.015625,0.0078125,-0.015625,0.0234375,-0.0078125,-0.0078125,0.0078125,-0.0078125,-0.0234375,-0.0234375,-0.0234375,0,-0.046875,0.0078125,0.03125,-0.0234375,-0.03125,-0.0078125,0.0078125,0,-0.0234375,-0.046875,-0.0390625,0.046875,0.0234375,-0.0078125,0,-0.015625,-0.0078125,-0.046875,0.0078125,-0.0546875,0,0.171875,0.03125,-0.0078125,0,-0.0078125,0.0078125,0.0078125,0.0078125,0.015625,0.0078125,0.0078125,0,-0.03125,-0.0234375,0.046875,-0.03125,-0.1015625,0.0703125,0.046875,-0.0390625,0,-0.0546875,0,-0.046875,-0.0078125,-0.0625,0.03125,0.046875,-0.0078125,-0.0234375,-0.015625,-0.0078125,-0.0234375,-0.1328125,-0.078125,-0.03125,0.09375,0.0234375,-0.015625,-0.0390625,-0.03125,-0.0390625,0.03125,-0.0234375,0,-0.0625,0.0390625,-0.0234375,-0.0078125,0.015625,-0.0234375,-0.015625,-0.046875,0.0234375,0.0390625,-0.0390625,0,-0.0078125,0.0078125,-0.0625,0.09375,0.03125,-0.0078125,0.0078125,-0.015625,0.0390625,0.0078125,-0.015625,0,-0.0703125,0.0390625,0.015625,0.03125,-0.0234375,0,-0.0078125,-0.0078125,0.0078125,-0.046875,-0.015625,-0.046875,-0.0234375,-0.0234375,-0.0234375,-0.015625,-0.015625,-0.0859375,0.046875,-0.0859375,-0.0546875,0.03125,0,-0.0390625,-0.015625,-0.0078125,-0.0390625,0.0390625,0.0390625,0.0078125,0.0078125,0.03125,0,0,-0.0078125,0,-0.0078125,0,-0.0234375,0.015625,-0.0078125,-0.015625,0.0078125,-0.015625,-0.015625,0,0,-0.015625,-0.0390625,-0.0078125,-0.015625,-0.0234375,-0.015625,0.03125,0.0390625,0.140625,-0.046875,0,0.0625,-0.015625,0,0.0078125,-0.0234375,0.0390625,0.03125,0.0234375,0.0625,-0.0625,0,-0.0390625,0.0078125,-0.015625,0.0703125,-0.015625,-0.0390625,-0.0390625,-0.0234375,0,-0.03125,-0.015625,-0.0625,0,-0.015625,0,-0.09375,0.015625,0.0078125,-0.0078125,0,-0.0546875,-0.0234375,-0.015625,-0.078125,0.015625,-0.0390625,-0.015625,-0.015625,-0.015625,-0.0234375,-0.09375,0.03125,-0.0234375,-0.0703125,0.015625,-0.0390625,-0.0234375,-0.015625,-0.0078125,0.0546875,-0.0859375,-0.015625,0.0390625,0.046875,0.0234375,-0.0078125,0.015625,-0.0390625,-0.0390625,-0.0234375,-0.0859375,0.1328125,-0.0078125,0.03125,0.0390625,0,0.0234375,-0.1328125,-0.015625,-0.0390625,-0.015625,-0.0546875,0,-0.0078125,-0.03125,-0.0234375,-0.03125,-0.03125,0.1015625,-0.046875,0.0625,-0.0078125,0.0078125,-0.0078125,0.046875,0.03125,0.0078125,0.03125,-0.03125,-0.078125,0.03125,0.03125,-0.0234375,0.0078125,-0.09375,0.0703125,0.0234375,-0.0625,-0.0546875,0.0390625,0,0.015625,0.0546875,-0.078125,-0.0546875,-0.015625,0.015625,-0.0078125,0,-0.015625,-0.015625,-0.0546875,0.0390625,0.1171875,-0.0078125,-0.0625,-0.046875,-0.03125,0.03125,0.125,-0.015625,-0.0234375,0,0.0078125,-0.0234375,-0.0078125,-0.0078125,-0.0078125,0.015625,-0.0078125,-0.015625,-0.015625,0,-0.0078125,-0.0078125,0,-0.09375,-0.09375,0,-0.0078125,-0.0078125,0,0.015625,0,-0.03125,-0.0703125,-0.03125,-0.015625,0.046875,-0.0078125,-0.015625,0.0234375,0,-0.0078125,-0.0390625,-0.015625,-0.0078125,-0.0390625,-0.109375,0.0078125,-0.0546875,0.03125,-0.0078125,0.0078125,0.015625,-0.015625,0,-0.015625,-0.0078125,0,0,-0.015625,-0.0234375,0.0234375,-0.0078125,0,-0.03125,-0.015625,-0.015625,-0.03125,-0.0078125,0.0625,0.078125,-0.03125,-0.03125,-0.0234375,0,0.0078125,0.0078125,0.015625,0.046875,0.0390625,-0.03125,-0.09375,0.03125,0.0078125,-0.03125,0.0234375,-0.015625,-0.078125,0.0078125,-0.0234375,0.0234375,0.0703125,0.015625,0.0234375,0.0078125,-0.0234375,-0.0234375,0.0859375,0,-0.0078125,-0.0078125,0,0,-0.0703125,0,0.0078125,0,-0.0078125,0,0.03125,-0.015625,-0.0078125,-0.0078125,0.0078125,0.0078125,0,0.0078125,0,0.0234375,-0.0078125,0.015625,-0.0078125,-0.015625,-0.015625,-0.0078125,0,0.015625,0.0078125,-0.03125,0.0390625,0.046875,0,0,0.0078125,0,0.046875,-0.0625,0.03125,0.0390625,-0.0078125,0.03125,-0.046875,-0.0390625,0.0078125,-0.046875,0.046875,0.0234375,-0.03125,-0.046875,0,-0.0078125,-0.015625,0,0.0078125,-0.015625,0.0078125,-0.0078125,0.015625,-0.0234375,-0.015625,0.015625,-0.03125,0,0,-0.03125,-0.0390625,-0.0234375,-0.015625,-0.03125,-0.0625,-0.015625,0.0625,-0.0234375,0.015625,0.109375,-0.03125,0,0.03125,-0.03125,-0.0234375,-0.046875,-0.0546875,0.03125,0.0625,0.0546875,-0.0078125,0.0390625,-0.125,-0.0078125,0.03125,-0.125,0,0.0234375,0.0859375,-0.0234375,0.03125,0.0078125,-0.015625,-0.0234375,-0.0234375,0.0078125,-0.046875,0.0078125,-0.0234375,0.046875,-0.0390625,0.0234375,-0.0234375,-0.078125,0.0234375,-0.015625,0.0234375,-0.015625,0.03125,-0.0546875,-0.0078125,0.0390625,0.1640625,-0.0234375,0.09375,-0.0625,-0.0078125,-0.015625,0.0390625,-0.015625,-0.03125,-0.0234375,-0.0078125,-0.046875,-0.0546875,-0.0078125,-0.046875,0.046875,-0.0234375,0.0234375,-0.0390625,-0.03125,0.03125,-0.0234375,0,0.046875,0.0234375,-0.015625,0.015625,-0.0625,0.0078125,-0.0703125,0.0859375,0.015625,0.0390625,-0.0625,0,-0.0703125,0.0390625,-0.0390625,-0.03125,-0.0390625,-0.0390625,-0.015625,-0.0078125,-0.0390625,-0.0390625,-0.109375,-0.0078125,0.015625,0.09375,-0.0234375,-0.0625,-0.0078125,-0.03125,0.0703125,0,-0.0078125,-0.0546875,-0.03125,-0.03125,0,0.0390625,-0.015625,-0.046875,-0.0546875,0.0078125,0.0078125,-0.0546875,-0.0078125,0.109375,0.1484375,-0.015625,-0.0390625,0.03125,0,-0.0390625,-0.0390625,0.015625,-0.0546875,0.0078125,0.078125,0.0078125,-0.0390625,-0.046875,-0.078125,-0.015625,0.0078125,0,0.0078125,0.0078125,-0.0078125,0,0.0078125,-0.015625,0,-0.046875,0.0390625,0.0078125,-0.0390625,-0.0703125,-0.0078125,0.0390625,-0.0703125,-0.0234375,0.0234375,-0.0234375,0.015625,0.0390625,-0.0390625,0.015625,0.0625,-0.0546875,0.0078125,0,-0.0234375,-0.0390625,0.015625,0,-0.0078125,-0.03125,0.0546875,0.015625,0,-0.0078125,0.0078125,0.0078125,0,0,0.0078125,-0.0078125,-0.0078125,0.015625,-0.0390625,-0.0234375,-0.0078125,0.03125,-0.0390625,-0.0234375,0.015625,0,-0.0859375,0.03125,0.03125,0.0859375,-0.0625,-0.015625,0.0078125,-0.078125,-0.015625,0.0625,-0.0234375,0.0234375,0.015625,-0.0078125,0.015625,-0.0625,0.0234375,-0.0234375,-0.0234375,0.0390625,0.03125,0.015625,-0.0390625,-0.0078125,0.046875,0.0078125,0.0078125,0,-0.015625,-0.0078125,-0.03125,-0.0234375,-0.0078125,0.015625,-0.0703125,0.015625,0.0078125,0.015625,0.015625,-0.0625,-0.03125,-0.0234375,0.03125,-0.03125,0.0234375,0,0.0078125,0.0234375,0,0,0,0.0078125,-0.0234375,-0.015625,0.0078125,-0.015625,-0.015625,-0.0234375,0.0234375,0,0.0546875,-0.03125,-0.015625,0.078125,-0.03125,-0.0078125,-0.078125,-0.0859375,0.0234375,0.0546875,-0.109375,-0.0078125,-0.03125,0.0078125,0.015625,0,0.09375,-0.03125,-0.109375,0.0078125,0.015625,-0.015625,0.0078125,0.015625,-0.015625,-0.0078125,-0.0078125,0,0,0,-0.046875,-0.03125,0.0078125,-0.015625,-0.0078125,-0.0078125,-0.015625,-0.015625,-0.0234375,0.015625,0,0.0078125,-0.015625,-0.0390625,-0.046875,0.1171875,-0.0703125,-0.015625,0.0078125,-0.03125,-0.03125,0.171875,-0.0546875,0.0078125,0.1640625,-0.0625,-0.0078125,0.0390625,0.0078125,0.0390625,-0.1015625,-0.015625,-0.03125,0.046875,0.03125,-0.0234375,0.0078125,-0.015625,0.0859375,-0.046875,-0.0078125,0,0.0078125,0.0390625,0.015625,0.0390625,0.0390625,-0.0390625,-0.0625,0.046875,-0.0390625,-0.0234375,-0.0546875,-0.0078125,-0.046875,-0.0390625,0.0078125,0.0390625,0.0234375,0,0.1015625,-0.09375,-0.0234375,0.0078125,0.0078125,-0.0234375,0.0625,0.0078125,-0.0234375,-0.0078125,0.015625,-0.0078125,-0.015625,0.09375,-0.0078125,-0.1171875,-0.0078125,-0.015625,-0.0390625,-0.0625,-0.046875,-0.0859375,0.03125,0.0234375,0.0078125,-0.078125,-0.015625,-0.046875,0.015625,0.015625,0.015625,0.015625,-0.0390625,-0.0546875,-0.046875,-0.0234375,0.125,-0.0078125,-0.0625,-0.03125,-0.03125,-0.0234375,-0.03125,-0.0625,0.0078125,0.1015625,0,0.0078125,-0.0625,0.046875,0.0078125,-0.078125,0,0.015625,0.0234375,-0.0078125,-0.0390625,0.0390625,0.0625,-0.015625,-0.0703125,-0.0078125,-0.015625,0,-0.03125,0.0078125,-0.0078125,0,0.0078125,0.09375,0.0234375,-0.03125,-0.046875,-0.0625,-0.0078125,-0.0390625,0.03125,0.1328125,-0.0078125,-0.0234375,0.0234375,0,-0.015625,-0.015625,0,0.0078125,0.0078125,-0.0078125,-0.0078125,0.015625,0,0.0078125,0,0.0234375,0.0390625,-0.0625,0.046875,0.0234375,-0.0078125,-0.015625,-0.015625,-0.0078125,-0.046875,0.046875,-0.015625,-0.046875,0.1015625,0.0234375,0,-0.015625,-0.03125,0.03125,-0.0625,-0.0078125,0.0078125,-0.0234375,0.0625,-0.0078125,0.0390625,0,-0.0078125,0.0078125,0,-0.015625,0.0078125,0,-0.015625,-0.0078125,-0.015625,-0.0078125,0.0703125,0,0.0078125,-0.03125,-0.03125,-0.0078125,0.0078125,0.0390625,-0.0390625,-0.0078125,-0.015625,-0.0625,-0.03125,0.078125,-0.0078125,0.015625,0,0.0078125,-0.0078125,0.015625,0.015625,0.015625,-0.03125,-0.0390625,-0.0546875,-0.046875,0.015625,-0.015625,0.0078125,0,-0.078125,0,-0.015625,-0.03125,-0.0390625,-0.03125,0,-0.0078125,-0.046875,0.0234375,0.0078125,-0.0078125,-0.0390625,0.03125,-0.0078125,0.015625,0.046875,-0.0078125,0,0.0390625,0,0.0234375,-0.015625,-0.0234375,0.0078125,-0.0546875,-0.015625,-0.0078125,-0.0078125,0.0078125,-0.0078125,-0.0078125,0.0390625,-0.015625,-0.0390625,-0.046875,0.0625,0.0234375,0,-0.0234375,0.03125,0.0078125,-0.078125,0.046875,-0.0078125,0.0078125,0.0234375,0,-0.0546875,-0.0078125,0.046875,0.03125,0,0.03125,0.0078125,-0.0703125,-0.03125,-0.015625,0.0234375,0,0,-0.0078125,0.0078125,0.015625,0.015625,0,0.0078125,0.0234375,-0.015625,-0.0078125,-0.015625,-0.0078125,-0.0390625,-0.03125,-0.0234375,0.0078125,-0.0078125,-0.03125,0.015625,0.0078125,-0.0234375,0.078125,-0.046875,0,-0.0234375,0.0078125,0.0078125,-0.03125,0.0859375,0.0390625,-0.0078125,0.0234375,-0.03125,0.0078125,-0.046875,0.015625,-0.0546875,0.0703125,-0.0390625,-0.109375,-0.1015625,0.03125,0.03125,0.0078125,0,-0.0625,-0.0078125,0.0078125,0.015625,0,-0.0078125,0.0390625,-0.015625,-0.0234375,0.0234375,-0.0078125,0.0078125,-0.0078125,-0.0234375,-0.015625,0,0,-0.0078125,0.0234375,0.015625,0.015625,-0.0703125,-0.015625,-0.046875,-0.015625,-0.0390625,-0.0625,0.0546875,-0.0078125,-0.0078125,-0.015625,0.0625,-0.0078125,0.0234375,-0.0234375,0,-0.0546875,-0.078125,0,0.0234375,0.0390625,0.0078125,0,0.046875,0,0.0078125,-0.03125,0.0234375,-0.03125,0,0.0078125,0.0234375,0.0234375,0.03125,0.0703125,-0.046875,-0.0078125,0.015625,-0.1015625,0.03125,-0.03125,0,0.0078125,-0.046875,-0.09375,-0.03125,0.015625,0,0.0078125,-0.046875,0.078125,0.0625,-0.015625,-0.046875,-0.03125,0.015625,0,-0.015625,-0.1015625,0.03125,0.0546875,-0.1015625,-0.0078125,-0.0078125,-0.0625,-0.015625,0,-0.015625,-0.015625,-0.0078125,0.0546875,0,-0.046875,-0.046875,-0.0078125,-0.03125,-0.046875,-0.015625,-0.0234375,0.0078125,0.0546875,-0.0390625,-0.0703125,0.0234375,0.0078125,0.0078125,0.0546875,0,-0.0078125,-0.0078125,-0.0078125,-0.0078125,-0.0078125,0,0,0,-0.0234375,0.0546875,0.09375,0.03125,-0.0234375,-0.109375,-0.0078125,0.0078125,-0.0078125,-0.015625,0.0078125,0.0078125,-0.015625,0.0546875,-0.078125,0.0078125,-0.0546875,0,0.046875,0.046875,-0.0234375,-0.03125,-0.0078125,-0.1328125,-0.078125,-0.03125,0.0078125,0.0078125,0.0078125,0.0234375,0,0.0078125,0,0,-0.0078125,-0.015625,-0.015625,0.0078125,-0.0703125,0.078125,0.0703125,-0.0078125,-0.015625,-0.1015625,-0.03125,-0.0390625,-0.0390625,-0.046875,-0.046875,-0.0625,-0.0078125,-0.015625,0.03125,0.1171875,-0.0078125,0.03125,0.03125,0.015625,-0.03125,-0.078125,-0.0234375,0.046875,0.0390625,-0.015625,-0.03125,-0.015625,0.046875,-0.0703125,-0.125,0.03125,0.0390625,0.1015625,0.0234375,0.0078125,-0.0234375,0,-0.0859375,-0.0234375,0.0078125,0.03125,-0.0625,0,0.0234375,-0.046875,-0.0078125,0.0234375,0.0703125,-0.015625,0.0078125,0.03125,-0.015625,0.0078125,0.015625,0.0078125,0,0.09375,-0.015625,0,0,0,-0.0078125,0.0703125,0.0234375,-0.0078125,-0.0546875,-0.046875,-0.03125,-0.046875,-0.015625,0.03125,-0.0703125,-0.03125,-0.015625,-0.0625,-0.0078125,0.0859375,0.0390625,0.0234375,0,-0.0546875,0.0078125,0.0078125,0,0.0078125,0,0.0625,-0.015625,-0.0078125,-0.0078125,-0.0078125,-0.0390625,-0.0078125,0.0078125,0.0078125,0.015625,-0.015625,0.03125,-0.0390625,0,-0.03125,0.0234375,0.0390625,-0.0546875,0.03125,0.0078125,-0.0546875,0.0234375,-0.015625,-0.046875,0.03125,-0.0078125,-0.0546875,0.0234375,-0.0078125,-0.015625,-0.0390625,-0.046875,0.03125,-0.078125,0,0.078125,0,0.0234375,-0.046875,0.125,0.0078125,-0.1171875,0,-0.0625,-0.046875,0.046875,-0.0234375,0.0546875,-0.1171875,-0.03125,-0.0234375,-0.0390625,-0.03125,0.046875,0.09375,0.015625,-0.046875,0.046875,-0.03125,0,-0.0234375,0.015625,0.046875,-0.0234375,0,0.0234375,0.0234375,-0.0078125,-0.0546875,-0.0234375,-0.0625,0.0234375,-0.0078125,0.0078125,0.0390625,-0.0703125,-0.03125,-0.015625,-0.0546875,0.0078125,0,0.125,0.0390625,-0.0546875,0,0,-0.03125,0.03125,-0.015625,0.03125,0.0546875,-0.0234375,-0.015625,0.125,-0.0078125,-0.0234375,-0.0546875,-0.0234375,0.0625,0.0625,-0.03125,0.015625,0.0234375,0.015625,-0.0546875,0.140625,0.0234375,-0.078125,0.0234375,0.0625,-0.03125,0.1171875,0.0078125,-0.046875,0.0234375,-0.0703125,-0.0234375,-0.1015625,0.03125,0.0234375,0.03125,0.03125,-0.015625,-0.1171875,-0.015625,0.046875,-0.125,0.0703125,-0.0390625,0.109375,-0.0078125,-0.125,-0.109375,0.0078125,0.0234375,-0.0546875,0.015625,0.0390625,-0.0625,0.0234375,-0.03125,0.0078125,-0.015625,-0.0390625,-0.0625,-0.0390625,-0.0625,-0.015625,-0.015625,0.0859375,0.09375,0.0078125,-0.078125,-0.046875,0,-0.015625,-0.0078125,-0.0078125,-0.0078125,0,-0.015625,0,0.0078125,0.015625,0.0546875,-0.0078125,-0.0078125,-0.0859375,-0.03125,-0.0078125,0.0234375,-0.046875,0.015625,0,-0.015625,0.015625,0.0625,-0.03125,-0.0390625,0.015625,-0.0078125,0.0078125,0,0.0078125,0.0234375,0.0703125,-0.0546875,-0.0078125,-0.03125,-0.03125,-0.0078125,-0.015625,0.0078125,-0.0078125,0,0.0078125,-0.0078125,0.0078125,0,-0.015625,0.0234375,0,0,0.03125,-0.078125,-0.015625,-0.046875,-0.046875,0.0234375,0.0546875,-0.0625,-0.0078125,-0.0859375,-0.0703125,0.0390625,0.0390625,0.015625,-0.03125,0.0625,-0.015625,0.015625,0.015625,-0.046875,0.0234375,0.0078125,-0.046875,-0.015625,-0.03125,0.0234375,0,-0.0078125,-0.0390625,-0.0078125,-0.0078125,-0.0078125,-0.0390625,0,0.015625,0,-0.046875,0,0.0078125,-0.0546875,-0.0859375,-0.015625,-0.0234375,0,-0.015625,-0.015625,0.0390625,-0.015625,-0.0078125,0,0.015625,0.0234375,-0.0078125,-0.015625,-0.0078125,0.015625,-0.0078125,-0.0078125,0.046875,0.0234375,0.0390625,0.03125,-0.0078125,-0.0390625,-0.0078125,-0.0234375,-0.0390625,-0.09375,-0.0390625,-0.015625,-0.046875,0.015625,0.078125,-0.0703125,-0.0234375,0,-0.0078125,0,0,-0.03125,-0.015625,-0.015625,0.0390625,-0.0234375,-0.0234375,0.1015625,0,-0.0078125,0,-0.0078125,0.0078125,0,-0.0078125,0,-0.015625,0.0390625,0,-0.0078125,-0.0078125,-0.046875,0.0234375,-0.0234375,0.015625,-0.0078125,0.015625,-0.0390625,-0.015625,-0.015625,-0.0234375,-0.0078125,0.0078125,-0.0546875,-0.0390625,-0.015625,-0.0078125,-0.0625,-0.03125,0.0625,0.0234375,-0.015625,-0.046875,-0.0859375,0.0078125,-0.078125,0.03125,-0.015625,-0.03125,0.1171875,-0.0390625,0,-0.0390625,0.0234375,-0.046875,-0.0390625,-0.0390625,0.0390625,-0.1015625,-0.0390625,0,0.1171875,-0.03125,-0.0390625,0.03125,-0.0234375,-0.0234375,0.0546875,-0.0390625,-0.0078125,-0.046875,0.0078125,-0.015625,-0.0078125,-0.0234375,-0.015625,0.0546875,-0.015625,-0.015625,-0.046875,-0.0078125,-0.0546875,-0.0078125,0.015625,-0.0625,-0.0078125,-0.0078125,0.03125,0,0.015625,-0.046875,0.046875,-0.046875,-0.109375,-0.0078125,-0.0234375,-0.0234375,0.0078125,0.0625,0.0625,-0.0234375,-0.0390625,0.0546875,0.015625,0.0078125,-0.046875,0.046875,0.0078125,-0.0078125,-0.1171875,-0.03125,-0.0078125,0.0703125,-0.0078125,-0.0234375,0.171875,0.0078125,-0.015625,0.0078125,-0.015625,-0.03125,0.015625,0,-0.03125,-0.046875,0.015625,0.0078125,-0.046875,-0.046875,-0.0703125,-0.109375,0,0.125,-0.1484375,-0.0078125,0.03125,0.046875,-0.015625,-0.078125,0.125,-0.0390625,-0.03125,-0.109375,0,-0.0546875,0.0390625,-0.0390625,0.0859375,-0.0234375,0.015625,-0.0078125,0,0.046875,-0.0234375,-0.0078125,0.0078125,-0.0234375,0.0078125,-0.015625,-0.0234375,0.046875,0.0078125,0.0078125,-0.0078125,-0.0078125,0.015625,-0.0078125,0,0,0.0078125,0.015625,-0.03125,0.015625,-0.015625,0,-0.015625,-0.046875,0.046875,0.0234375,0.0703125,-0.03125,-0.0234375,-0.0390625,-0.0390625,0.1171875,-0.0546875,-0.078125,0.0390625,-0.0703125,0.078125,-0.0078125,-0.0390625,-0.0078125,-0.0234375,-0.015625,0.0234375,-0.03125,-0.0078125,0.0078125,-0.015625,0,0.0078125,-0.0078125,0.0078125,-0.0078125,0.0078125,0.1015625,0.0234375,0.0234375,0.0625,-0.0234375,-0.0390625,-0.046875,-0.015625,-0.0546875,0.0703125,0,-0.03125,0.03125,-0.015625,0.03125,-0.03125,0.0703125,-0.0078125,0.0078125,-0.046875,0.015625,-0.1015625,-0.09375,0.0390625,0.0546875,-0.0625,-0.0234375,0.015625,0.0234375,-0.0078125,-0.03125,-0.03125,0.0078125,0.0625,0.1015625,0.046875,0.046875,0.0703125,0.0546875,0.046875,-0.03125,-0.0390625,-0.015625,0.0390625,-0.03125,-0.0078125,-0.03125,0.03125,0.0390625,0.0703125,0.03125,-0.0234375,-0.0390625,-0.015625,-0.046875,-0.0546875,-0.03125,0.015625,0.046875,-0.0078125,-0.015625,0.015625,0.0078125,0.0078125,-0.015625,-0.0234375,0.0625,-0.015625,-0.0078125,-0.0390625,-0.046875,-0.0234375,0.0625,0.0859375,-0.0078125,-0.0703125,-0.046875,-0.0703125,0,0.0390625,0.0625,0.015625,0.03125,0.0859375,-0.0078125,-0.0703125,-0.0625,0,0,0.015625,0.0078125,0,0.0078125,0.015625,0.015625,0.0078125,0.0078125,-0.0078125,-0.0078125,0.0234375,-0.0078125,-0.0546875,0.0390625,-0.03125,0.046875,-0.0390625,0.0078125,0.03125,0.0078125,-0.0546875,-0.0390625,-0.0703125,-0.0625,-0.03125,0.0625,-0.046875,-0.0234375,-0.0078125,0.0546875,0,-0.0859375,0.015625,-0.0234375,-0.0234375,0.03125,-0.0859375,0.03125,0.0859375,0.0390625,0.0078125,-0.0078125,-0.0703125,-0.0234375,0.015625,0.0078125,-0.046875,0.0078125,-0.09375,-0.0078125,0.0390625,-0.0703125,0.0078125,0.046875,0.0703125,-0.0234375,-0.015625,0.015625,0.0234375,-0.0625,-0.015625,-0.015625,-0.0390625,0.0078125,-0.0859375,0.0625,0.09375,-0.078125,-0.03125,-0.046875,-0.046875,0.0234375,-0.0703125,0.0078125,0.0234375,-0.03125,-0.015625,0,-0.0234375,-0.0390625,-0.0078125,-0.03125,-0.0703125,-0.078125,0.0234375,-0.046875,-0.1015625,0,0,0.0078125,0.046875,-0.03125,-0.0625,-0.03125,0,-0.015625,0.0859375,-0.0859375,-0.046875,-0.0234375,-0.046875,0.0078125,0.03125,-0.015625,-0.0703125,-0.046875,-0.03125,-0.015625,0.0234375,0,0.078125,0,-0.03125,0.1015625,0,-0.0078125,0.0234375,-0.0546875,0.0546875,-0.0078125,0.015625,0.0859375,-0.0234375,-0.0234375,-0.0390625,-0.0078125,0,0.0390625,-0.03125,0.0390625,0.0078125,0.03125,-0.09375,-0.0234375,0.03125,0,-0.078125,-0.0078125,0.046875,0.125,-0.0625,0.015625,0.015625,0.0078125,0.046875,0.0234375,-0.0078125,0.015625,-0.015625,0,0.0625,-0.0703125,-0.0703125,0,-0.0078125,-0.0078125,0.0078125,0.015625,-0.015625,-0.015625,-0.015625,-0.0078125,-0.015625,0,-0.0390625,-0.046875,-0.09375,-0.109375,0.015625,0.0546875,0.0078125,-0.015625,0.015625,-0.078125,-0.03125,-0.015625,-0.015625,-0.0234375,-0.046875,-0.0390625,-0.0234375,-0.03125,-0.015625,-0.015625,0.015625,-0.03125,-0.015625,0.125,-0.03125,-0.0234375,0.0078125,-0.0078125,0,0,0.0078125,-0.0078125,0.0078125,0,0.0078125,-0.046875,-0.09375,-0.03125,-0.078125,0.03125,-0.0078125,-0.09375,0.125,0,-0.109375,0.0390625,-0.0078125,0.0078125,0,0.015625,-0.0859375,0,0,0.03125,-0.0078125,-0.0078125,0.1015625,-0.0859375,-0.0390625,0.0859375,-0.078125,-0.0390625,0.046875,-0.0234375,0.015625,-0.0234375,0.0234375,0.0078125,0.0078125,0.015625,0,0,0.0390625,-0.0390625,0.0234375,-0.015625,0.0078125,0,-0.0546875,-0.0078125,-0.0703125,-0.0234375,0.015625,0,0.0078125,-0.0078125,-0.03125,-0.0546875,-0.0234375,0,-0.0234375,0.0078125,-0.0390625,-0.015625,-0.0078125,-0.0390625,0.0234375,0,0.0625,-0.0078125,0,0.0390625,0.015625,-0.03125,0.0078125,-0.015625,-0.0078125,0.0625,-0.0546875,-0.03125,0.0234375,0.0625,0.015625,-0.109375,0,-0.0390625,-0.015625,-0.0546875,-0.0078125,-0.0859375,-0.03125,-0.0546875,0.0625,0,-0.03125,-0.0078125,-0.0234375,0,0.0078125,-0.0078125,-0.0078125,0.03125,0.0078125,0,-0.046875,-0.0546875,0,0.0234375,-0.015625,-0.0078125,0.0234375,0.0625,0.0078125,-0.0703125,-0.046875,-0.015625,0.0625,-0.0390625,-0.0234375,-0.0234375,0.0390625,-0.0234375,0,0.015625,-0.03125,-0.03125,-0.1015625,-0.03125,-0.0234375,-0.0625,-0.03125,0,-0.109375,-0.0078125,-0.0078125,-0.03125,0.0234375,-0.046875,0.1015625,0.015625,-0.03125,-0.0546875,-0.015625,-0.03125,0.0078125,0.0234375,0.125,-0.0234375,-0.03125,-0.0078125,-0.03125,-0.0390625,0.0625,-0.0390625,0.0234375,0.0234375,-0.0390625,-0.0078125,-0.046875,0.0546875,-0.03125,0.0859375,-0.015625,-0.078125,-0.03125,-0.03125,-0.0234375,-0.0625,-0.0625,-0.015625,0.03125,0.0390625,0.0078125,0.0234375,0.015625,0.0234375,-0.0078125,0.0625,-0.015625,0,-0.0546875,0.03125,0,0.03125,0,0.0234375,-0.0078125,0,-0.0625,-0.0234375,-0.015625,0.0234375,-0.03125,-0.0546875,0.0703125,-0.0078125,-0.046875,0.078125,0.0390625,-0.0625,-0.09375,-0.0546875,0.03125,0.046875,-0.0234375,-0.0078125,-0.0390625,-0.0390625,-0.0078125,0.078125,-0.0078125,0.0234375,-0.0078125,0.0078125,0,-0.0390625,0,-0.0234375,-0.03125,0,-0.0234375,-0.03125,0.0546875,-0.0234375,-0.03125,-0.0546875,-0.046875,0.015625,0.0625,-0.03125,-0.03125,0.09375,0.015625,0.046875,-0.0390625,-0.015625,-0.0078125,-0.0625,-0.015625};


outputs = '{0.125,0.1875,0.3125,0.125,0.125,0.1875,0.3125,0.125,0.125,0.25,0.125,0.0625,0.1875,0.1875,0.1875,0,0,0,0,0,0,0.0625,0.125,0,0,0,0.0625,0.3125,0.25,0.5,0.3125,0.0625,0.375,0.0625,0,0.0625,0,0,0,0.0625,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0.125,0,0.0625,0.4375,0.125,0.125,0,0,0,0,0,0,0,0.0625,0.0625,0,0,0,0,0,0,0,0,0,0,0.125,0.0625,0,0,0,0,0,0,0.4375,0.1875,0.25,0,0,0,0.1875,0,0,0.1875,0.0625,0.125,0,0,0.25,0,0,0,0.4375,0,0.375,0.1875,0.125,0.125,0.3125,0.0625,0.1875,0.375,0.1875,0.25,0,0,0,0,0.3125,0.1875,0,0.25,0.25,0.25,0.4375,0.5,0.375,0.1875,0.1875,0.1875,0,0,0.125,0.0625,0.0625,0.0625,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0.5625,0.125,0.375,0.1875,0.1875,0.25,0.125,0.0625,0.25,0,0,0,0.25,0,0.0625,0.125,0,0.1875,0,0,0,0,0,0,0,0.125,0,0.3125,0.125,0.3125,0.3125,0,0.3125,0.5,0.0625,0.3125,0.125,0.125,0.3125,0,0,0.1875,0.5,0.0625,0.3125,0,0,0,0,0,0,0,0,0,0,0,0,0,0.0625,0,0,0,0,0,0.1875,0.3125,0,0,0,0,0.125,0,0.375,0.1875,0.25,0.1875,0,0.1875,0,0,0,0.125,0,0.0625,0,0.0625,0,0,0,0,0.125,0.1875,0.125,0.125,0.125,0.0625,0,0.0625,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0.0625,0,0,0.0625,0,0.4375,0.4375,0.5,0.5,0.0625,0.25,0,0,0,0,0,0,0,0,0,0.0625,0,0,0.125,0.125,0.0625,0.0625,0.0625,0.1875,0,0,0,0,0,0,0,0.1875,0,0.0625,0.125,0.1875,0.0625,0,0,0,0,0.0625,0,0,0,0,0,0,0,0,0,0,0,0,0.1875,0.1875,0.0625,0.0625,0.0625,0,0,0,0,0.375,0.25,0.875,0.125,0,0.375,0,0,0,0,0,0,0,0,0,0.0625,0.1875,0.25,0.3125,0.3125,0.5,0.125,0.375,0.5,0,0.5,0.4375,0,0,0,0,0,0,0,0.125,0,0,0.3125,0.375,0,0,0.1875,0.375,0.0625,0.0625,0.375,0.5,0.375,0.25,0.1875,0.375,0,0.0625,0.0625,0,0,0.1875,0,0,0,0,0,0,0.3125,0.4375,0.1875,0.1875,0.1875,0.375,0,0,0,0.3125,0.125,0.125,0.0625,0,0,0.125,0.25,0,0.4375,0.5,0.5,0,0.25,0.4375,0,0,0,0.5625,0.125,0,0.0625,0.125,0.125,0.3125,0.375,0.3125,0.375,0.125,0.25,0.1875,0,0.0625,0,0.0625,0,0.1875,0.375,0.125,0.125,0.125,0.1875,0.1875,0.25,0.25,0,0,0,0,0.25,0,0.1875,0.375,0.3125,0.1875,0.25,0.3125,0.0625,0.0625,0.375,0.3125,0,0.1875,0,0,0,0,0,0,0,0.3125,0.125,0,0.125,0.0625,0.0625,0.375,0.25,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0.0625,0,0,0,0,0.125,0,0,0,0.1875,0.3125,0,0,0.1875,0,0,0,0,0.125,0.0625,0.0625,0,0.0625,0.3125,0.125,0.375,0.0625,0.1875,0.3125,0,0.0625,0,0,0,0.375,0,0,0.0625,0,0.0625,0,0,0,0,0,0.0625,0,0,0.375,0.1875,0.0625,0.0625,0,0,0,0.0625,0.125,0,0.0625,0.0625,0,0.1875,0,0,0,0,0,0,0,0,0,0.125,0,0,0,0,0,0.6875,0.125,0.0625,0.4375,0,0.0625,0.625,0.0625,0.25,0,0,0,0,0,0,0,0.0625,0.1875,0,0,0,0,0.25,0.125,0.125,0.125,0.25,0.0625,0.125,0.1875,0,0.0625,0.1875,0,0,0.0625,0.125,0.0625,0,0,0,0,0.3125,0,0,0,0,0,0,0,0,0,0.0625,0.125,0,0,0.0625,0.0625,0,0.0625,0.3125,0.0625,0.3125,0.6875,0.125,0.5625,0.3125,0.0625,0.3125,0,0.0625,0,0.125,0.0625,0.25,0,0,0.0625,0,0,0,0.1875,0,0,0.0625,0.0625,0.0625,0.4375,0.375,0.4375,0,0,0,0.0625,0.0625,0.0625,0,0,0,0.3125,0.125,0.3125,0.1875,0.0625,0.125,0.125,0,0.125,0.5625,0.3125,0.375,0.4375,0.125,0.375,0.4375,0.3125,0.5,0.4375,0.25,0.375,0.3125,0,0.1875,0,0,0,0,0,0.125,0,0,0.0625,0,0,0,0,0.125,0,0,0.25,0.1875,0.4375,0.1875,0.5,0.4375,0,0.625,0.5625,0.0625,0.375,0.6875,0.1875,0.375,0,0,0,0,0,0,0,0,0,0,0,0.5625,0.0625,0.1875,0.4375,0,0.1875,0.125,0.375,0.375,0.6875,0,0.0625,0.25,0.125,0.125,0.125,0.6875,0.4375,0.75,0.5625,0,0.5,0.375,0.0625,0.125,0,0,0,0,0,0,0.25,0.3125,0.125,0,0,0,0,0,0,0,0,0,0.0625,0.1875,0.5625,0,0,0,0,0,0,0.1875,0.0625,0.3125,0.0625,0,0.125,0,0,0,0.3125,0.375,0.8125,0.4375,0,0.5,0,0,0,0.125,0.0625,0,0.0625,0.1875,0,0.3125,0.25,0.25,0.125,0.125,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0.0625,0,0.0625,0.125,0,0,0,0,0,0,0,0,0,0,0,0,0.125,0,0,0,0.25,0,0,0,0,0,0,0.125,0,0,0.0625,0.1875,0,0.125,0.1875,0.25,0,0,0,0,0,0,0,0,0,0.3125,0.4375,0.375,0.25,0.125,0.5625,0.375,0.125,0.4375,0.3125,0.1875,0,0.1875,0.125,0,0.5,0.0625,0.125,0.8125,0.5625,0.8125,1.25,0.1875,0.6875,0.0625,0,0,0.125,0,0,0.125,0,0,0.125,0,0,0,0.1875,0.375,0,0,0.25,0,0.1875,0.25,0.125,0,0,0.0625,0.125,0.0625,0.1875,0,0,0,0,0,0,0,0,0,0.125,0.0625,0,0,0,0,0,0,0.75,0.125,0.5,0,0.0625,0.0625,0,0,0,0,0,0,0.375,0,0.25,0.1875,0,0,0.75,0.375,0.5,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0.0625,0.0625,0.125,0,0,0,0,0,0,0,0,0,0.0625,0,0,0,0.0625,0,0.1875,0.1875,0.0625,0,0,0,0,0.0625,0.0625,0.125,0.25,0.4375,0.1875,0.0625,0,0.125,0,0,0,0,0,0.1875,0.1875,0.5625,0,0,0,0.3125,0.125,0,0,0.125,0,0.0625,0,0,0.125,0.125,0,0,0,0,0,0,0,0.1875,0.125,0.25,0.375,0.125,0.6875,0.375,0,0.125,0.3125,0.125,0,0.3125,0,0.1875,0.125,0.0625,0,0,0,0,0,0,0,0,0,0,0,0,0,0.125,0.0625,0,0,0,0,0.0625,0.1875,0.1875,0.125,0.1875,0.125,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0.1875,0.1875,0.1875,0,0,0.125,0.4375,0.1875,0.5,0,0,0,0,0.0625,0.125,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0.5,0.25,0.375,0.5,0.375,0.75,0.25,0.0625,0.75,0,0,0,0.1875,0,0,0.4375,0,0,0.3125,0,0,0,0,0.25,0,0,0,0.4375,0,0,0.375,0.125,0.0625,0,0,0,0,0,0,0,0,0,0.0625,0,0,0.1875,0,0,0,0,0,0,0,0.125,0.375,0,0,0,0.375,0,0.9375,1.4375,0.1875,0,0.3125,0,0,0,0,0,0.4375,0.875,0,0.5,0.5,0.4375,0.25,0.25,0,0.625,0,0.1875,0.1875,0,0,0,0,0,0,0,0.4375,0.0625,0.375,0.0625,0,0,0.5625,0,0.3125,0.25,0,0.125,0.125,0.375,0.5,0,0,0.3125,0.0625,0,0.5,0,0,0,0.5625,0.125,0.125,0.125,0.0625,0,0.125,0,0.6875,0,0,0,0.5625,0,0.1875,0,0,0,0,0,0,0,0,0.125,0,0,0,0,0,0,0.1875,1.125,0.25,0,0,0.0625,0,0,0,0,0,0.1875,0,0.3125,0,0.3125,1.375,0,0,0,0,0.3125,0,0,0.375,0,0,0,0,0,0.125,0.0625,0,0,0.1875,0,0,0,0,0,0,0,0.1875,0.25,0,0,0,0,0,0,0,0,0.3125,0,0.25,0.1875,0.1875,0,0,0,0,0,0,0,0.0625,0,0,0.0625,0.25,0.125,0.3125,0.625,0,0,0.375,0,0,0,0,0,0.125,0.25,0,0.1875,0.3125,0.1875,0.5,0.4375,0,0.75,0.5625,0,0,0.75,0.125,0.0625,0,0,0,0,0.125,0,0,0.875,0,0,0,0,0,0.0625,0,0.25,0.25,0,0,0,0,0.125,0,0.125,0.625,0,0.3125,1.0,0,0,0.1875,0,0,0,0,0.1875,0,0.125,0.75,0,0,0,0.375,0.0625,0.5,0.375,0,0.1875,0,0,0.0625,0,0,0,0,0,0.375,0,0,0,0,0,0,0,0.375,0.125,0,0,0,0,0,0,0.5625,0,0,0.375,0,0.0625,0,0,0,0,0.5,0,0,0,0,0,0,0,0.0625,0,0,0.1875,0,0.0625,0.3125,0,0,0,0,0,0,0.6875,0,0,0,0,0.3125,0.9375,1.5,0,0,0.1875,0.6875,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0.125,0,0.1875,0.0625,0,0,0,0,0,0.6875,0.3125,0,0,0,0,0.5,0.875,0.4375,0.3125,0.5,0,0,0.1875,0.6875,0.125,0.6875,0,0.25,0.5625,0.6875,0.1875,0.625,0.125,0,0.1875,0,0.125,0,0,0,0,0,0,0,0,0,0,0,1.125,0,0,0.75,0,0,0,0,0,0.0625,0,0,0,0,0,0,0,0,0.3125,0,0,0.0625,0,0,0,0,0,0.25,0,0,0,0,0,0,0,0.25,0.1875,0,0.375,0.8125,0.4375,0,0.25,0.0625,0,0,0,0,0,0,0.1875,0,0.25,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0.125,0.125,0,0.5625,0.0625,0,0,0,0,0,0.375,0.0625,0.5,0,0.1875,0,0,0,0,0.4375,0,0,0,0,0,0,0,0,0,0,0.875,0,0,0,0.375,0,0,0.1875,0.0625,0.0625,0.0625,0.125,0.25,0.75,0.25,0,0,0,0,0,0,0,0.4375,0.6875,0.625,0.6875,0.75,0,0,0,0,0,0,0.1875,0,0,0.375,0.75,0.1875,0,0.1875,0,0,0,0,0,0,0,0,0,0.125,0,0,0.125,0,0,0.0625,0.0625,0.9375,0,0,0.8125,0,0,0.4375,0,0.0625,0,0,0.8125,0,0,0.3125,0.25,0,0,0,0,0,0,0,0.25,0.25,0,0,0,0,0.5625,0,0.5,0.75,0,0.5625,0,0,0,0,0.0625,0,0,0,0,0.6875,0,0,0.1875,0,0,0,0.375,0,0.1875,0.4375,0.25,0,0,0,0,0.25,0,0.25,1.0625,0.1875,0.75,1.4375,0.5,0,0,0,0,0.1875,0.0625,0,0,0,0.1875,0.125,0.125,0,0,0,0,0,0.0625,0,0,0,0.125,0,0,0,0,0.125,0,0,0.0625,0,0,0,0,0,0,0.375,0,0,0.3125,1.3125,0.375,0,1.0,0,0,0.6875,0,0,0,0,0.0625,0,0,0.1875,0,0.125,0,0,0,0,0,0,0.0625,0.3125,0,0.125,0,0,0.5,0.8125,0.9375,0.8125,0.1875,0.8125,0.5,0.5,0.8125,0,0,0,0.8125,0,0.4375,0,0,0,0,0,0.125,0,0.5625,0.6875,0,0.3125,0,0,0,0.125,0,0.0625,0.3125,0.25,0.4375,0.5,0,0,0,0.1875,0,0.25,0,0,0,0.1875,0.1875,0,0,0.4375,0,0.375,0,0,0,0,0,0,0,0,0,0,0,0.75,0,0.4375,0.3125,0,0.125,0,0,0,0,0,0,0,0,0,0,0,0,0.125,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1.0,0.3125,0.75,0.9375,0,1.1875,1.1875,1.125,0.9375,0,0,0,0,1.4375,1.0625,0,0.0625,0.5,0.1875,0.125,0,0.0625,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0.5,0.625,0.25,1.0,0.5625,0,0.0625,0.25,0,0,0,0,0,0,0,0,0.5625,0.3125,0,0,0.1875,0,0,0,0,0,0,0,0,0,0.375,0,0.0625,0.25,0.4375,0.8125,0.9375,0.75,0.5625,0.125,0.375,0,0,0,0,0.8125,0,0,1.0625,0,0,0.9375,0,0,0,0.0625,0,0,0.1875,0.25,0,0,0.25,0,0,0,0,0,0,0.0625,0,0.4375,0,0.5,0.5625,0,0.8125,0.3125,0.125,0.25,0,0,0,0,0.9375,0,0,0,0,0.6875,0,0.6875,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0.25,0,0.375,0.75,0,0.4375,0,0.75,0,0.4375,0.875,0.5625,0,0,0.0625,0,0.0625,0.75,0,0,0,0.0625,0.1875,0,0,0,0,0.75,1.125,0.6875,0,0,0,0.125,0.3125,0,0.0625,0.0625,0,0.0625,0,0.125,0,0,0,0.4375,0,0.3125,0,0,0,0.4375,0.3125,1.0625,0,0,0.8125,0.5,0.0625,0.75,0.25,0.5,0.3125,0,0,0,0.125,0,0.25,0.1875,0,0,0.5625,0,0,0,0.8125,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0.125,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0.1875,0,0,0.4375,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0.25,0,0,0.125,0,0,0,0,0,0,0,0,0.5,0.25,0.4375,0,0.5625,0.625,0.375,1.3125,0.125,0.5625,0.6875,0.25,0,0,0,0.375,0.0625,0.125,0.375,0.1875,0.5625,0,0,0,0.5,0,0.8125,0.5,0.0625,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0.4375,0.3125,0.0625,0.625};
        clk <= 0;

        counter <= 0;

        rst = 1'b1;
        for(int i = 0; i < 9; i++)begin
            PE_inputs[i] = 8'd0;
            PE_weights[i] = 8'd0;
        end
        #120;
        rst = 0;
        #40;
        bias3x3 <= 0;

        val = -8'd128;
        index = -8;
        for(int i = 0; i < 256; i++)begin
            lookup_input[index] = new[1];
            lookup_input[index] = '{val};
            index = index + 0.0625;
            val = val + 8'd1;
        end

        val = -8'd128;
        index = -8;
        for(int i = 0; i < 256; i++)begin
            lookup_output[index] = new[1];
            lookup_output[index] = '{val};
            index = index + 0.0625;
            val = val + 8'd1;
        end

        val = -8'd128;
        index = -1;
        for(int i = 0; i < 256; i++)begin
            lookup_weight[index] = new[1];
            lookup_weight[index] = '{val};
            index = index + 0.0078125;
            val = val + 8'd1;
        end

        // PE_weights[0] = 8'd4;
        // PE_inputs[0] = 8'd7;
        // #40;

        // rst <= 1'b1;
        // #40;
        // rst<=1'b0;
        // #40;

        for(int i = 0; i < 9; i++)begin
            PE_inputs[i] = 8'd0;
            PE_weights[i] = 8'd0;
        end
        #40;

			#20;

        for(int i =0; i < 32; i++)begin 
            for(int j = 0; j < 256; j++)begin//for loop for first convolution
                for(int k = 0; k < 9; k++)begin
                    PE_inputs[k] = lookup_input[inputs[j*9+k]][0];
                    PE_weights[k] = lookup_weight[weight_s[i*256+j]][0];
                end
                #40;
                counter <= counter + 1;
            end
            for(int w = 0; w < 9; w++)begin
                PE_weights[w] = lookup_weight[bias_s[i]][0];
                PE_inputs[w] = lookup_input[1][0];
            end
            #40;
            counter <= counter + 1;
            for(int k = 0; k < 9; k++)begin
//                output_s[i*9 + k] = new[1];
                output_s[i*9 + k] = PE_outputs[k];
            end
            rst <= 1'b1;
            for(int i = 0; i < 9; i++)begin
                PE_inputs[i] = 8'd0;
                PE_weights[i] = 8'd0;
            end
            #40;
            rst <= 1'b0;
            #40;
        end
			
			#40;
        //have to modify the first layer outputs to feed into other layers since clipping is different

        for(int i = 0; i < 128; i++)begin
            for(int j = 0; j < 32; j++)begin//for loop for the 1x1 expand
                for(int k = 0; k < 9; k++)begin
                    PE_inputs[k] = output_s[j*9+(8-k)];
                    PE_weights[k] = lookup_weight[weight_1x1[i*32+j]][0];
                end
                #40;
                counter <= counter + 1;    
            end
            for(int w = 0; w < 9; w++)begin
                PE_weights[w] = lookup_weight[bias_1x1[i]][0];
                PE_inputs[w] = lookup_input[1][0];
            end
            #40;
            counter <= counter + 1;
            for(int k = 0; k < 9; k++)begin
//                output_[i*9 + k] = new[1];
                output_[i*9 + k] = PE_outputs[k];
            end
            rst <= 1'b1;
            for(int i = 0; i < 9; i++)begin
                PE_inputs[i] = 8'd0;
                PE_weights[i] = 8'd0;
            end
            #40;
            rst <= 1'b0;
            #40;
        end

        for(int i = 0; i < 128; i++)begin//for loop for the 3x3 expand
            for(int j = 0; j < 9; j++)begin
                for(int k = 0; k < 32; k++)begin
                    for(int w = 0; w < 9; w++)begin
                        PE_weights[w] = lookup_weight[weight_3x3[i*32*9+k*9+w]][0];
                    end
                    if(j==0)begin
                        PE_inputs[0] = lookup_input[0][0];
                        PE_inputs[1] = lookup_input[0][0];
                        PE_inputs[2] = lookup_input[0][0];
                        PE_inputs[3] = lookup_input[0][0];
                        PE_inputs[4] = output_s[k*9+8];
                        PE_inputs[5] = output_s[k*9+7];
                        PE_inputs[6] = lookup_input[0][0];
                        PE_inputs[7] = output_s[k*9+5];
                        PE_inputs[8] = output_s[k*9+4];
                    end
                    else if(j==1)begin
                        PE_inputs[0] = lookup_input[0][0];
                        PE_inputs[1] = lookup_input[0][0];
                        PE_inputs[2] = lookup_input[0][0];
                        PE_inputs[3] = output_s[k*9+8];
                        PE_inputs[4] = output_s[k*9+7];
                        PE_inputs[5] = output_s[k*9+6];
                        PE_inputs[6] = output_s[k*9+5];
                        PE_inputs[7] = output_s[k*9+4];
                        PE_inputs[8] = output_s[k*9+3];
                    end
                    else if(j==2)begin
                        PE_inputs[0] = lookup_input[0][0];
                        PE_inputs[1] = lookup_input[0][0];
                        PE_inputs[2] = lookup_input[0][0];
                        PE_inputs[3] = output_s[k*9+7];
                        PE_inputs[4] = output_s[k*9+6];
                        PE_inputs[5] = lookup_input[0][0];
                        PE_inputs[6] = output_s[k*9+4];
                        PE_inputs[7] = output_s[k*9+3];
                        PE_inputs[8] = lookup_input[0][0];
                    end
                    else if(j==3)begin
                        PE_inputs[0] = lookup_input[0][0];
                        PE_inputs[1] = output_s[k*9+8];
                        PE_inputs[2] = output_s[k*9+7];
                        PE_inputs[3] = lookup_input[0][0];
                        PE_inputs[4] = output_s[k*9+5];
                        PE_inputs[5] = output_s[k*9+4];
                        PE_inputs[6] = lookup_input[0][0];
                        PE_inputs[7] = output_s[k*9+2];
                        PE_inputs[8] = output_s[k*9+1];
                    end
                    else if(j==4)begin
                        PE_inputs[0] = output_s[k*9+8];
                        PE_inputs[1] = output_s[k*9+7];
                        PE_inputs[2] = output_s[k*9+6];
                        PE_inputs[3] = output_s[k*9+5];
                        PE_inputs[4] = output_s[k*9+4];
                        PE_inputs[5] = output_s[k*9+3];
                        PE_inputs[6] = output_s[k*9+2];
                        PE_inputs[7] = output_s[k*9+1];
                        PE_inputs[8] = output_s[k*9];
                    end
                    else if(j==5)begin
                        PE_inputs[0] = output_s[k*9+7];
                        PE_inputs[1] = output_s[k*9+6];
                        PE_inputs[2] = lookup_input[0][0];
                        PE_inputs[3] = output_s[k*9+4];
                        PE_inputs[4] = output_s[k*9+5];
                        PE_inputs[5] = lookup_input[0][0];
                        PE_inputs[6] = output_s[k*9+1];
                        PE_inputs[7] = output_s[k*9];
                        PE_inputs[8] = lookup_input[0][0];
                    end
                    else if(j==6)begin
                        PE_inputs[0] = lookup_input[0][0];
                        PE_inputs[1] = output_s[k*9+5];
                        PE_inputs[2] = output_s[k*9+4];
                        PE_inputs[3] = lookup_input[0][0];
                        PE_inputs[4] = output_s[k*9+2];
                        PE_inputs[5] = output_s[k*9+1];
                        PE_inputs[6] = lookup_input[0][0];
                        PE_inputs[7] = lookup_input[0][0];
                        PE_inputs[8] = lookup_input[0][0];
                    end
                    else if(j==7)begin
                        PE_inputs[0] = output_s[k*9+5];
                        PE_inputs[1] = output_s[k*9+4];
                        PE_inputs[2] = output_s[k*9+3];
                        PE_inputs[3] = output_s[k*9+2];
                        PE_inputs[4] = output_s[k*9+1];
                        PE_inputs[5] = output_s[k*9];
                        PE_inputs[6] = lookup_input[0][0];
                        PE_inputs[7] = lookup_input[0][0];
                        PE_inputs[8] = lookup_input[0][0];
                    end
                    else if(j==8)begin
                        PE_inputs[0] = output_s[k*9+4];
                        PE_inputs[1] = output_s[k*9+3];
                        PE_inputs[2] = lookup_input[0][0];
                        PE_inputs[3] = output_s[k*9+1];
                        PE_inputs[4] = output_s[k*9];
                        PE_inputs[5] = lookup_input[0][0];
                        PE_inputs[6] = lookup_input[0][0];
                        PE_inputs[7] = lookup_input[0][0];
                        PE_inputs[8] = lookup_input[0][0];
                    end
                    #40;
                    counter <= counter + 1;
                end
                bias3x3 = lookup_weight[bias_3x3[i]][0];
                #40;
                bias3x3 = 8'b0;
                counter <= counter + 1;
//                output_3x3[i*9+j] = new[1];
                output_3x3[i*9+j] = out_3x3; 
                rst <= 1'b1;
                for(int i = 0; i < 9; i++)begin
                    PE_inputs[i] = 8'd0;
                    PE_weights[i] = 8'd0;
                end
                #40;
                rst <= 1'b0;
                #40;
            end
        end
		  
		  #40;

        //compare the ideal outputs 
        for(int i = 0; i < 1152; i++)begin
            if(output_[i] != lookup_output[outputs[i]][0])begin
                   $error("Output wrong at index %d. DUT:0x%h, BASELINE:0x%h", i,
                   output_[i], lookup_output[outputs[i]][0]); 
            end
        end
        for(int i = 0; i < 1152; i++)begin
            if(output_3x3[i] != lookup_output[outputs[i+1152]][0])begin
                   $error("Output wrong at index %d. DUT:0x%h, BASELINE:0x%h", i+1152,
						 output_3x3[i], lookup_output[outputs[i+1152]][0]); 
            end
        end
		$finish;
    end
	 
endmodule
