package arrays;

inputs = [0.125,0.1875,0.3125,0.125,0.125,0.1875,0.3125,0.125,0.125,0.25,0.125,0.0625,0.1875,0.1875,0.1875,0.0,0.0,0.0,0.0,0.0,0.0,0.0625,0.125,0.0,0.0,0.0,0.0625,0.3125,0.25,0.5,0.3125,0.0625,0.375,0.0625,0.0,0.0625,0.0,0.0,0.0,0.0625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.125,0.0,0.0625,0.4375,0.125,0.125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0625,0.0625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.125,0.0625,0.0,0.0,0.0,0.0,0.0,0.0,0.4375,0.1875,0.25,0.0,0.0,0.0,0.1875,0.0,0.0,0.1875,0.0625,0.125,0.0,0.0,0.25,0.0,0.0,0.0,0.4375,0.0,0.375,0.1875,0.125,0.125,0.3125,0.0625,0.1875,0.375,0.1875,0.25,0.0,0.0,0.0,0.0,0.3125,0.1875,0.0,0.25,0.25,0.25,0.4375,0.5,0.375,0.1875,0.1875,0.1875,0.0,0.0,0.125,0.0625,0.0625,0.0625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.5625,0.125,0.375,0.1875,0.1875,0.25,0.125,0.0625,0.25,0.0,0.0,0.0,0.25,0.0,0.0625,0.125,0.0,0.1875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.125,0.0,0.3125,0.125,0.3125,0.3125,0.0,0.3125,0.5,0.0625,0.3125,0.125,0.125,0.3125,0.0,0.0,0.1875,0.5,0.0625,0.3125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0625,0.0,0.0,0.0,0.0,0.0,0.1875,0.3125,0.0,0.0,0.0,0.0,0.125,0.0,0.375,0.1875,0.25,0.1875,0.0,0.1875,0.0,0.0,0.0,0.125,0.0,0.0625,0.0,0.0625,0.0,0.0,0.0,0.0,0.125,0.1875,0.125,0.125,0.125,0.0625,0.0,0.0625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0625,0.0,0.0,0.0625,0.0,0.4375,0.4375,0.5,0.5,0.0625,0.25,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0625,0.0,0.0,0.125,0.125,0.0625,0.0625,0.0625,0.1875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1875,0.0,0.0625,0.125,0.1875,0.0625,0.0,0.0,0.0,0.0,0.0625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1875,0.1875,0.0625,0.0625,0.0625,0.0,0.0,0.0,0.0,0.375,0.25,0.875,0.125,0.0,0.375,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0625,0.1875,0.25,0.3125,0.3125,0.5,0.125,0.375,0.5,0.0,0.5,0.4375,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.125,0.0,0.0,0.3125,0.375,0.0,0.0,0.1875,0.375,0.0625,0.0625,0.375,0.5,0.375,0.25,0.1875,0.375,0.0,0.0625,0.0625,0.0,0.0,0.1875,0.0,0.0,0.0,0.0,0.0,0.0,0.3125,0.4375,0.1875,0.1875,0.1875,0.375,0.0,0.0,0.0,0.3125,0.125,0.125,0.0625,0.0,0.0,0.125,0.25,0.0,0.4375,0.5,0.5,0.0,0.25,0.4375,0.0,0.0,0.0,0.5625,0.125,0.0,0.0625,0.125,0.125,0.3125,0.375,0.3125,0.375,0.125,0.25,0.1875,0.0,0.0625,0.0,0.0625,0.0,0.1875,0.375,0.125,0.125,0.125,0.1875,0.1875,0.25,0.25,0.0,0.0,0.0,0.0,0.25,0.0,0.1875,0.375,0.3125,0.1875,0.25,0.3125,0.0625,0.0625,0.375,0.3125,0.0,0.1875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.3125,0.125,0.0,0.125,0.0625,0.0625,0.375,0.25,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0625,0.0,0.0,0.0,0.0,0.125,0.0,0.0,0.0,0.1875,0.3125,0.0,0.0,0.1875,0.0,0.0,0.0,0.0,0.125,0.0625,0.0625,0.0,0.0625,0.3125,0.125,0.375,0.0625,0.1875,0.3125,0.0,0.0625,0.0,0.0,0.0,0.375,0.0,0.0,0.0625,0.0,0.0625,0.0,0.0,0.0,0.0,0.0,0.0625,0.0,0.0,0.375,0.1875,0.0625,0.0625,0.0,0.0,0.0,0.0625,0.125,0.0,0.0625,0.0625,0.0,0.1875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.125,0.0,0.0,0.0,0.0,0.0,0.6875,0.125,0.0625,0.4375,0.0,0.0625,0.625,0.0625,0.25,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0625,0.1875,0.0,0.0,0.0,0.0,0.25,0.125,0.125,0.125,0.25,0.0625,0.125,0.1875,0.0,0.0625,0.1875,0.0,0.0,0.0625,0.125,0.0625,0.0,0.0,0.0,0.0,0.3125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0625,0.125,0.0,0.0,0.0625,0.0625,0.0,0.0625,0.3125,0.0625,0.3125,0.6875,0.125,0.5625,0.3125,0.0625,0.3125,0.0,0.0625,0.0,0.125,0.0625,0.25,0.0,0.0,0.0625,0.0,0.0,0.0,0.1875,0.0,0.0,0.0625,0.0625,0.0625,0.4375,0.375,0.4375,0.0,0.0,0.0,0.0625,0.0625,0.0625,0.0,0.0,0.0,0.3125,0.125,0.3125,0.1875,0.0625,0.125,0.125,0.0,0.125,0.5625,0.3125,0.375,0.4375,0.125,0.375,0.4375,0.3125,0.5,0.4375,0.25,0.375,0.3125,0.0,0.1875,0.0,0.0,0.0,0.0,0.0,0.125,0.0,0.0,0.0625,0.0,0.0,0.0,0.0,0.125,0.0,0.0,0.25,0.1875,0.4375,0.1875,0.5,0.4375,0.0,0.625,0.5625,0.0625,0.375,0.6875,0.1875,0.375,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.5625,0.0625,0.1875,0.4375,0.0,0.1875,0.125,0.375,0.375,0.6875,0.0,0.0625,0.25,0.125,0.125,0.125,0.6875,0.4375,0.75,0.5625,0.0,0.5,0.375,0.0625,0.125,0.0,0.0,0.0,0.0,0.0,0.0,0.25,0.3125,0.125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0625,0.1875,0.5625,0.0,0.0,0.0,0.0,0.0,0.0,0.1875,0.0625,0.3125,0.0625,0.0,0.125,0.0,0.0,0.0,0.3125,0.375,0.8125,0.4375,0.0,0.5,0.0,0.0,0.0,0.125,0.0625,0.0,0.0625,0.1875,0.0,0.3125,0.25,0.25,0.125,0.125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0625,0.0,0.0625,0.125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.125,0.0,0.0,0.0,0.25,0.0,0.0,0.0,0.0,0.0,0.0,0.125,0.0,0.0,0.0625,0.1875,0.0,0.125,0.1875,0.25,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.3125,0.4375,0.375,0.25,0.125,0.5625,0.375,0.125,0.4375,0.3125,0.1875,0.0,0.1875,0.125,0.0,0.5,0.0625,0.125,0.8125,0.5625,0.8125,1.25,0.1875,0.6875,0.0625,0.0,0.0,0.125,0.0,0.0,0.125,0.0,0.0,0.125,0.0,0.0,0.0,0.1875,0.375,0.0,0.0,0.25,0.0,0.1875,0.25,0.125,0.0,0.0,0.0625,0.125,0.0625,0.1875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.125,0.0625,0.0,0.0,0.0,0.0,0.0,0.0,0.75,0.125,0.5,0.0,0.0625,0.0625,0.0,0.0,0.0,0.0,0.0,0.0,0.375,0.0,0.25,0.1875,0.0,0.0,0.75,0.375,0.5,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0625,0.0625,0.125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0625,0.0,0.0,0.0,0.0625,0.0,0.1875,0.1875,0.0625,0.0,0.0,0.0,0.0,0.0625,0.0625,0.125,0.25,0.4375,0.1875,0.0625,0.0,0.125,0.0,0.0,0.0,0.0,0.0,0.1875,0.1875,0.5625,0.0,0.0,0.0,0.3125,0.125,0.0,0.0,0.125,0.0,0.0625,0.0,0.0,0.125,0.125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1875,0.125,0.25,0.375,0.125,0.6875,0.375,0.0,0.125,0.3125,0.125,0.0,0.3125,0.0,0.1875,0.125,0.0625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.125,0.0625,0.0,0.0,0.0,0.0,0.0625,0.1875,0.1875,0.125,0.1875,0.125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1875,0.1875,0.1875,0.0,0.0,0.125,0.4375,0.1875,0.5,0.0,0.0,0.0,0.0,0.0625,0.125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.5,0.25,0.375,0.5,0.375,0.75,0.25,0.0625,0.75,0.0,0.0,0.0,0.1875,0.0,0.0,0.4375,0.0,0.0,0.3125,0.0,0.0,0.0,0.0,0.25,0.0,0.0,0.0,0.4375,0.0,0.0,0.375,0.125,0.0625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0625,0.0,0.0,0.1875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.125,0.375,0.0,0.0,0.0,0.375,0.0,0.9375,1.4375,0.1875,0.0,0.3125,0.0,0.0,0.0,0.0,0.0,0.4375,0.875,0.0,0.5,0.5,0.4375,0.25,0.25,0.0,0.625,0.0,0.1875,0.1875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.4375,0.0625,0.375,0.0625,0.0,0.0,0.5625,0.0,0.3125,0.25,0.0,0.125,0.125,0.375,0.5,0.0,0.0,0.3125,0.0625,0.0,0.5,0.0,0.0,0.0,0.5625,0.125,0.125,0.125,0.0625,0.0,0.125,0.0,0.6875,0.0,0.0,0.0,0.5625,0.0,0.1875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.125,0.0,0.0,0.0,0.0,0.0,0.0,0.1875,1.125,0.25,0.0,0.0,0.0625,0.0,0.0,0.0,0.0,0.0,0.1875,0.0,0.3125,0.0,0.3125,1.375,0.0,0.0,0.0,0.0,0.3125,0.0,0.0,0.375,0.0,0.0,0.0,0.0,0.0,0.125,0.0625,0.0,0.0,0.1875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1875,0.25,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.3125,0.0,0.25,0.1875,0.1875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0625,0.0,0.0,0.0625,0.25,0.125,0.3125,0.625,0.0,0.0,0.375,0.0,0.0,0.0,0.0,0.0,0.125,0.25,0.0,0.1875,0.3125,0.1875,0.5,0.4375,0.0,0.75,0.5625,0.0,0.0,0.75,0.125,0.0625,0.0,0.0,0.0,0.0,0.125,0.0,0.0,0.875,0.0,0.0,0.0,0.0,0.0,0.0625,0.0,0.25,0.25,0.0,0.0,0.0,0.0,0.125,0.0,0.125,0.625,0.0,0.3125,1.0,0.0,0.0,0.1875,0.0,0.0,0.0,0.0,0.1875,0.0,0.125,0.75,0.0,0.0,0.0,0.375,0.0625,0.5,0.375,0.0,0.1875,0.0,0.0,0.0625,0.0,0.0,0.0,0.0,0.0,0.375,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.375,0.125,0.0,0.0,0.0,0.0,0.0,0.0,0.5625,0.0,0.0,0.375,0.0,0.0625,0.0,0.0,0.0,0.0,0.5,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0625,0.0,0.0,0.1875,0.0,0.0625,0.3125,0.0,0.0,0.0,0.0,0.0,0.0,0.6875,0.0,0.0,0.0,0.0,0.3125,0.9375,1.5,0.0,0.0,0.1875,0.6875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.125,0.0,0.1875,0.0625,0.0,0.0,0.0,0.0,0.0,0.6875,0.3125,0.0,0.0,0.0,0.0,0.5,0.875,0.4375,0.3125,0.5,0.0,0.0,0.1875,0.6875,0.125,0.6875,0.0,0.25,0.5625,0.6875,0.1875,0.625,0.125,0.0,0.1875,0.0,0.125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.125,0.0,0.0,0.75,0.0,0.0,0.0,0.0,0.0,0.0625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.3125,0.0,0.0,0.0625,0.0,0.0,0.0,0.0,0.0,0.25,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.25,0.1875,0.0,0.375,0.8125,0.4375,0.0,0.25,0.0625,0.0,0.0,0.0,0.0,0.0,0.0,0.1875,0.0,0.25,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.125,0.125,0.0,0.5625,0.0625,0.0,0.0,0.0,0.0,0.0,0.375,0.0625,0.5,0.0,0.1875,0.0,0.0,0.0,0.0,0.4375,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.875,0.0,0.0,0.0,0.375,0.0,0.0,0.1875,0.0625,0.0625,0.0625,0.125,0.25,0.75,0.25,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.4375,0.6875,0.625,0.6875,0.75,0.0,0.0,0.0,0.0,0.0,0.0,0.1875,0.0,0.0,0.375,0.75,0.1875,0.0,0.1875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.125,0.0,0.0,0.125,0.0,0.0,0.0625,0.0625,0.9375,0.0,0.0,0.8125,0.0,0.0,0.4375,0.0,0.0625,0.0,0.0,0.8125,0.0,0.0,0.3125,0.25,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.25,0.25,0.0,0.0,0.0,0.0,0.5625,0.0,0.5,0.75,0.0,0.5625,0.0,0.0,0.0,0.0,0.0625,0.0,0.0,0.0,0.0,0.6875,0.0,0.0,0.1875,0.0,0.0,0.0,0.375,0.0,0.1875,0.4375,0.25,0.0,0.0,0.0,0.0,0.25,0.0,0.25,1.0625,0.1875,0.75,1.4375,0.5,0.0,0.0,0.0,0.0,0.1875,0.0625,0.0,0.0,0.0,0.1875,0.125,0.125,0.0,0.0,0.0,0.0,0.0,0.0625,0.0,0.0,0.0,0.125,0.0,0.0,0.0,0.0,0.125,0.0,0.0,0.0625,0.0,0.0,0.0,0.0,0.0,0.0,0.375,0.0,0.0,0.3125,1.3125,0.375,0.0,1.0,0.0,0.0,0.6875,0.0,0.0,0.0,0.0,0.0625,0.0,0.0,0.1875,0.0,0.125,0.0,0.0,0.0,0.0,0.0,0.0,0.0625,0.3125,0.0,0.125,0.0,0.0,0.5,0.8125,0.9375,0.8125,0.1875,0.8125,0.5,0.5,0.8125,0.0,0.0,0.0,0.8125,0.0,0.4375,0.0,0.0,0.0,0.0,0.0,0.125,0.0,0.5625,0.6875,0.0,0.3125,0.0,0.0,0.0,0.125,0.0,0.0625,0.3125,0.25,0.4375,0.5,0.0,0.0,0.0,0.1875,0.0,0.25,0.0,0.0,0.0,0.1875,0.1875,0.0,0.0,0.4375,0.0,0.375,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.75,0.0,0.4375,0.3125,0.0,0.125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.0,0.3125,0.75,0.9375,0.0,1.1875,1.1875,1.125,0.9375,0.0,0.0,0.0,0.0,1.4375,1.0625,0.0,0.0625,0.5,0.1875,0.125,0.0,0.0625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.5,0.625,0.25,1.0,0.5625,0.0,0.0625,0.25,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.5625,0.3125,0.0,0.0,0.1875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.375,0.0,0.0625,0.25,0.4375,0.8125,0.9375,0.75,0.5625,0.125,0.375,0.0,0.0,0.0,0.0,0.8125,0.0,0.0,1.0625,0.0,0.0,0.9375,0.0,0.0,0.0,0.0625,0.0,0.0,0.1875,0.25,0.0,0.0,0.25,0.0,0.0,0.0,0.0,0.0,0.0,0.0625,0.0,0.4375,0.0,0.5,0.5625,0.0,0.8125,0.3125,0.125,0.25,0.0,0.0,0.0,0.0,0.9375,0.0,0.0,0.0,0.0,0.6875,0.0,0.6875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.25,0.0,0.375,0.75,0.0,0.4375,0.0,0.75,0.0,0.4375,0.875,0.5625,0.0,0.0,0.0625,0.0,0.0625,0.75,0.0,0.0,0.0,0.0625,0.1875,0.0,0.0,0.0,0.0,0.75,1.125,0.6875,0.0,0.0,0.0,0.125,0.3125,0.0,0.0625,0.0625,0.0,0.0625,0.0,0.125,0.0,0.0,0.0,0.4375,0.0,0.3125,0.0,0.0,0.0,0.4375,0.3125,1.0625,0.0,0.0,0.8125,0.5,0.0625,0.75,0.25,0.5,0.3125,0.0,0.0,0.0,0.125,0.0,0.25,0.1875,0.0,0.0,0.5625,0.0,0.0,0.0,0.8125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1875,0.0,0.0,0.4375,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.25,0.0,0.0,0.125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.5,0.25,0.4375,0.0,0.5625,0.625,0.375,1.3125,0.125,0.5625,0.6875,0.25,0.0,0.0,0.0,0.375,0.0625,0.125,0.375,0.1875,0.5625,0.0,0.0,0.0,0.5,0.0,0.8125,0.5,0.0625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.4375,0.3125,0.0625,0.625];

bias_s = [0.03125,0.0078125,-0.1015625,0.0,0.21875,-0.015625,0.09375,0.3359375,0.15625,0.0,0.109375,0.1328125,0.0234375,-0.078125,-0.046875,0.0859375,0.03125,-0.0390625,0.078125,0.1328125,0.03125,0.03125,0.203125,-0.0625,0.09375,0.0,-0.0234375,0.0703125,-0.0703125,0.0078125,0.21875,0.0];

bias_1x1 = [-0.015625,-0.015625,-0.046875,-0.015625,-0.0,-0.0703125,0.0234375,-0.015625,-0.046875,0.015625,-0.03125,-0.0234375,-0.0390625,-0.015625,-0.078125,0.015625,-0.015625,-0.015625,0.03125,-0.0078125,0.0078125,-0.015625,-0.0390625,0.0078125,0.03125,-0.015625,-0.0234375,0.0234375,-0.015625,-0.0390625,-0.0,-0.0078125,-0.03125,-0.03125,-0.0390625,-0.0234375,-0.0390625,-0.0078125,-0.015625,-0.0078125,-0.0234375,-0.0078125,-0.0078125,-0.046875,0.0078125,-0.03125,-0.015625,-0.0,-0.015625,-0.0234375,-0.03125,-0.0390625,0.0,-0.03125,-0.0,-0.0234375,-0.0234375,-0.0078125,-0.0,-0.015625,-0.0625,-0.0,-0.015625,-0.0390625,-0.0234375,-0.0078125,-0.0234375,-0.015625,0.0,-0.0078125,-0.03125,0.0234375,-0.015625,-0.09375,0.0078125,0.015625,-0.015625,-0.03125,-0.015625,-0.0546875,-0.0234375,-0.0390625,0.015625,-0.015625,-0.0,-0.0078125,-0.0234375,0.0078125,-0.0078125,-0.0,-0.03125,-0.1015625,-0.015625,-0.0234375,-0.0234375,-0.0,-0.03125,-0.046875,-0.0078125,-0.03125,-0.015625,0.0,-0.015625,-0.046875,-0.046875,-0.0546875,-0.0546875,-0.0546875,-0.015625,-0.0234375,-0.0234375,-0.0078125,-0.03125,-0.015625,-0.015625,0.0078125,-0.03125,-0.0078125,-0.0859375,-0.015625,-0.0390625,-0.0234375,-0.0078125,-0.0234375,-0.0234375,0.015625,-0.046875,-0.0390625];

bias_3x3 = [-0.015625,-0.046875,-0.0078125,0.0390625,-0.0,-0.09375,-0.015625,-0.0546875,-0.015625,-0.09375,-0.0859375,-0.0234375,-0.015625,-0.0078125,-0.0390625,-0.03125,0.0234375,-0.0546875,-0.046875,-0.0234375,0.046875,-0.046875,-0.0390625,-0.0390625,-0.078125,0.0234375,-0.0703125,-0.046875,-0.1171875,-0.0546875,-0.0078125,0.0078125,-0.0390625,-0.0546875,-0.015625,-0.0078125,0.0,-0.0546875,-0.0546875,-0.046875,-0.0,-0.0078125,-0.0234375,-0.0546875,-0.03125,-0.03125,0.0390625,-0.015625,-0.03125,-0.0234375,0.0078125,-0.0234375,-0.078125,-0.0625,-0.015625,-0.0234375,-0.0546875,-0.0703125,-0.0234375,-0.0546875,0.0078125,-0.0234375,-0.0234375,-0.0,-0.0546875,0.015625,0.0234375,0.0078125,-0.0078125,0.0,0.046875,-0.046875,-0.0234375,-0.09375,-0.0703125,0.03125,-0.0,-0.046875,-0.125,0.0078125,-0.1171875,0.0,0.0234375,-0.0234375,0.0078125,-0.03125,-0.0546875,0.0234375,-0.0703125,-0.0703125,-0.046875,-0.0625,0.0078125,-0.0390625,-0.0546875,-0.015625,0.0078125,0.03125,0.0,-0.0078125,-0.03125,-0.0390625,-0.0625,0.0390625,-0.015625,-0.0078125,-0.015625,-0.03125,0.0,0.0390625,0.078125,-0.1171875,-0.0625,-0.0625,-0.0546875,-0.0625,-0.0,-0.046875,-0.046875,-0.03125,0.0234375,-0.015625,0.015625,0.0078125,0.015625,0.0234375,-0.015625,0.015625];

weight_s = [-0.03125,0.0078125,0.03125,-0.015625,0.0,-0.0078125,0.0703125,-0.0234375,-0.03125,-0.0859375,0.0546875,-0.109375,-0.03125,0.0234375,0.03125,0.015625,0.0078125,-0.0390625,0.0,-0.0,-0.0625,-0.0859375,0.046875,0.0,0.0390625,-0.0390625,-0.015625,0.03125,-0.0078125,-0.015625,-0.0390625,0.03125,0.0,0.0234375,0.03125,-0.015625,0.0078125,-0.0,-0.0703125,0.0078125,-0.0234375,-0.03125,0.0078125,0.0859375,-0.0234375,-0.0078125,-0.078125,-0.109375,0.0234375,0.015625,0.046875,-0.046875,0.03125,0.0859375,-0.0078125,-0.0078125,0.0234375,0.015625,-0.0234375,0.0625,-0.1015625,-0.046875,-0.0,-0.0390625,-0.0390625,-0.0390625,0.1171875,0.015625,-0.046875,0.0859375,-0.0390625,0.0078125,-0.015625,-0.078125,-0.0234375,-0.015625,-0.0546875,0.0078125,-0.0,-0.0078125,-0.0234375,-0.0078125,0.1328125,0.0078125,-0.0234375,-0.0234375,-0.0078125,-0.0234375,-0.015625,-0.0,-0.03125,-0.0234375,-0.0078125,0.0,0.0078125,0.015625,-0.078125,-0.0078125,-0.0625,-0.0703125,0.0546875,0.0390625,0.0546875,-0.0390625,-0.0078125,0.0078125,0.0703125,-0.046875,-0.0078125,0.046875,0.046875,-0.0390625,0.0078125,0.015625,-0.0390625,0.015625,0.0390625,0.0703125,-0.046875,0.015625,-0.0390625,-0.03125,0.0,-0.03125,-0.0703125,-0.0234375,-0.046875,-0.015625,-0.0703125,-0.1015625,-0.046875,-0.1171875,0.0859375,0.171875,-0.03125,-0.0625,-0.0,0.1171875,0.125,-0.015625,-0.2265625,-0.015625,-0.09375,-0.1015625,0.109375,-0.0390625,-0.15625,0.03125,-0.0234375,0.015625,0.109375,-0.046875,-0.1796875,-0.0703125,0.0703125,-0.03125,0.0390625,0.0703125,-0.0390625,-0.1484375,-0.109375,-0.2109375,0.0234375,0.078125,-0.0234375,0.296875,0.0703125,-0.0390625,0.0625,-0.0703125,0.0625,0.03125,0.0625,-0.09375,0.140625,-0.1328125,0.0859375,0.140625,0.078125,0.03125,0.015625,-0.0625,-0.0,0.078125,0.0703125,-0.109375,0.0859375,-0.078125,0.1171875,-0.0703125,-0.0625,-0.015625,-0.0546875,-0.0390625,-0.0703125,0.03125,-0.046875,-0.0234375,0.0234375,0.2421875,-0.0078125,-0.140625,-0.1640625,0.0390625,0.0078125,0.046875,-0.015625,0.0,-0.03125,0.046875,-0.09375,-0.0234375,0.0234375,0.0390625,0.0234375,-0.0078125,-0.046875,0.0234375,-0.015625,0.1328125,-0.0390625,-0.0234375,0.1171875,-0.0390625,0.109375,0.03125,0.203125,0.140625,-0.0625,-0.1328125,-0.046875,-0.0,-0.0625,-0.0234375,0.140625,0.0703125,-0.078125,0.0,0.109375,0.0,-0.0078125,-0.0546875,0.1171875,0.03125,-0.1015625,0.1015625,-0.0390625,-0.109375,-0.0625,0.1328125,0.0859375,0.1640625,0.015625,-0.0234375,-0.078125,0.046875,0.0234375,0.0234375,0.0078125,-0.015625,-0.015625,-0.0078125,-0.0234375,0.03125,0.0234375,0.0625,-0.0078125,-0.015625,0.0078125,-0.015625,-0.015625,0.0078125,-0.0078125,-0.0078125,-0.0,0.015625,0.0,0.015625,-0.0078125,0.0078125,-0.0,0.0078125,-0.0078125,-0.0078125,0.0078125,-0.015625,0.0078125,-0.015625,-0.0,0.0,0.0234375,0.03125,-0.0234375,-0.0234375,0.0234375,-0.0390625,0.0234375,-0.0,0.0078125,-0.015625,0.015625,0.0078125,0.0,0.0234375,0.015625,0.015625,0.015625,0.015625,0.0078125,0.015625,0.015625,0.0,0.03125,0.0234375,0.015625,-0.0234375,0.03125,0.015625,0.0078125,0.015625,-0.0078125,0.0078125,0.015625,0.0078125,0.015625,0.0234375,-0.015625,0.0078125,-0.015625,0.015625,-0.015625,-0.0078125,-0.015625,0.0078125,0.0,0.015625,0.015625,0.015625,-0.015625,0.0,0.03125,0.015625,-0.0078125,-0.0234375,-0.0234375,-0.0234375,0.015625,0.0234375,-0.0078125,0.0078125,0.0078125,-0.015625,0.0390625,0.0,0.0078125,0.015625,-0.0390625,0.0078125,-0.015625,0.0078125,-0.0,-0.0078125,-0.015625,-0.015625,-0.0,0.015625,-0.0078125,-0.0078125,-0.0078125,0.015625,0.0,0.015625,-0.0,0.0,-0.0,-0.0078125,0.0078125,-0.0,0.015625,0.0,0.015625,0.015625,0.0,-0.0078125,0.0,-0.0078125,-0.0078125,0.0,0.015625,-0.0,0.015625,-0.0078125,-0.0234375,-0.0078125,-0.0078125,-0.0234375,-0.0078125,0.0,0.0,0.0078125,-0.0234375,0.015625,0.015625,0.0078125,-0.0,0.0078125,-0.0234375,-0.0234375,-0.0234375,-0.03125,0.015625,-0.0078125,-0.015625,0.03125,-0.0234375,-0.03125,-0.0078125,-0.0,0.0078125,-0.0,-0.0,0.0078125,-0.03125,0.03125,0.0234375,0.015625,0.015625,0.0234375,0.0,0.0234375,0.015625,-0.015625,0.0078125,-0.0078125,-0.0,-0.015625,0.0078125,-0.0078125,0.015625,0.03125,0.0,-0.015625,-0.015625,-0.015625,-0.0078125,-0.015625,-0.0078125,0.015625,-0.03125,0.0078125,-0.0234375,0.0234375,0.0078125,0.015625,-0.0078125,-0.015625,0.015625,0.0078125,-0.0078125,-0.015625,-0.0234375,-0.0078125,-0.0234375,0.0234375,0.0078125,-0.0078125,0.015625,0.0234375,0.0234375,0.0078125,0.03125,-0.0078125,-0.015625,-0.0078125,-0.0625,0.015625,0.0,0.015625,-0.0078125,0.0234375,-0.0078125,0.0,0.0078125,0.015625,-0.0234375,-0.0234375,-0.0078125,0.046875,-0.0078125,-0.015625,-0.03125,-0.015625,-0.015625,-0.0,0.0078125,-0.0,-0.0078125,-0.0078125,0.03125,-0.0,0.0078125,-0.0,-0.0,0.0,-0.0234375,-0.0078125,-0.0390625,-0.0234375,-0.015625,-0.0078125,0.015625,-0.0078125,0.0859375,0.078125,0.0078125,0.046875,-0.0234375,-0.0078125,-0.0,0.1171875,-0.0078125,-0.1328125,-0.0625,-0.0078125,0.0,-0.046875,0.0078125,-0.0,-0.0,0.0703125,-0.0078125,0.046875,0.015625,0.0390625,0.109375,-0.03125,-0.0390625,0.1015625,0.0234375,-0.0390625,0.0078125,0.015625,0.015625,-0.0078125,-0.015625,0.1171875,0.0546875,-0.0,-0.0078125,0.1328125,-0.0546875,0.0390625,-0.03125,0.03125,-0.03125,0.078125,0.046875,0.0234375,0.1640625,0.03125,0.015625,0.0546875,-0.1015625,0.046875,-0.0078125,0.0390625,0.0390625,0.0078125,0.0546875,-0.0546875,0.0390625,0.0078125,-0.0,0.0078125,-0.0234375,-0.015625,0.015625,0.0078125,-0.0546875,0.0234375,-0.046875,-0.0078125,-0.0234375,0.046875,0.0703125,-0.03125,0.03125,-0.03125,-0.0078125,0.046875,0.0625,-0.0390625,0.0546875,0.0,0.15625,0.0703125,0.09375,-0.03125,-0.0078125,0.046875,0.03125,0.140625,-0.0078125,-0.015625,0.0234375,0.015625,0.015625,0.125,0.0,0.03125,0.0625,-0.046875,0.0390625,-0.0078125,0.0703125,0.0234375,-0.0078125,-0.0546875,0.0234375,-0.0234375,-0.0078125,-0.078125,0.0078125,-0.015625,-0.015625,0.0390625,0.0625,0.0234375,0.0234375,0.0625,0.0078125,-0.0078125,-0.0,0.09375,-0.0,-0.03125,0.0546875,-0.046875,-0.0625,0.0703125,0.078125,0.0859375,-0.0390625,-0.0859375,0.1171875,0.0703125,-0.0234375,0.0390625,-0.046875,-0.0390625,-0.046875,-0.0546875,-0.125,-0.0390625,-0.0703125,-0.046875,0.0078125,0.0078125,-0.03125,0.015625,-0.0859375,0.0390625,0.125,0.078125,0.09375,0.0234375,0.0390625,-0.0078125,0.140625,-0.0390625,-0.09375,-0.09375,-0.109375,-0.1796875,0.046875,0.0078125,0.015625,-0.015625,0.109375,0.078125,-0.0703125,0.0546875,-0.0703125,-0.0234375,0.0390625,-0.0546875,0.1640625,-0.03125,-0.0625,0.0390625,-0.109375,-0.046875,0.0390625,0.046875,0.015625,-0.0625,-0.0390625,0.0390625,-0.0703125,0.015625,0.0,0.0390625,-0.0,0.09375,0.0234375,-0.0546875,-0.0546875,-0.1015625,0.015625,0.015625,0.0625,0.078125,-0.0234375,0.0390625,-0.03125,-0.0703125,-0.046875,-0.0390625,0.0078125,-0.1640625,-0.0234375,-0.0390625,-0.1015625,0.0078125,-0.1015625,-0.0859375,-0.0625,0.03125,0.140625,0.1015625,0.015625,0.203125,0.09375,-0.078125,0.1171875,0.046875,-0.171875,0.0703125,0.0078125,0.2421875,-0.015625,-0.109375,-0.046875,-0.0625,0.0546875,0.0546875,-0.0703125,-0.0078125,0.1015625,-0.046875,-0.0,0.046875,0.0625,0.09375,-0.09375,-0.0078125,0.0546875,0.0234375,-0.0234375,-0.140625,0.015625,0.015625,-0.03125,-0.0234375,-0.015625,0.0859375,0.109375,-0.0234375,0.0390625,0.03125,-0.0546875,-0.0,0.0078125,0.0078125,-0.0390625,-0.09375,-0.0234375,-0.03125,0.015625,-0.0390625,-0.0078125,0.0859375,0.015625,-0.015625,0.0078125,-0.0234375,0.015625,0.0078125,-0.0625,-0.03125,-0.03125,-0.0,0.0625,0.0546875,0.0078125,0.046875,0.0234375,-0.0390625,0.0625,0.046875,-0.0234375,0.0234375,-0.0234375,-0.0546875,-0.0,0.0078125,-0.0390625,0.1640625,-0.03125,0.015625,0.0859375,0.0546875,0.015625,0.0703125,0.0546875,0.03125,0.0234375,-0.0078125,-0.0390625,-0.0078125,0.1015625,-0.09375,-0.015625,-0.0390625,0.03125,-0.0078125,0.0859375,0.0625,-0.0078125,0.046875,-0.015625,-0.0390625,-0.078125,-0.0546875,-0.0546875,-0.0,-0.0390625,-0.015625,-0.0,0.109375,-0.0390625,0.0625,0.046875,-0.03125,0.0390625,0.03125,0.03125,-0.0234375,-0.0,0.0,0.0625,0.0078125,0.0234375,0.0703125,-0.0078125,-0.0078125,0.0234375,-0.015625,-0.0390625,-0.0234375,-0.0078125,0.0,0.03125,0.0078125,-0.03125,-0.015625,0.0078125,-0.03125,0.03125,-0.0390625,0.0390625,-0.0234375,-0.03125,-0.046875,-0.0078125,-0.015625,-0.0078125,-0.015625,-0.03125,-0.0,0.015625,0.0234375,0.0078125,-0.0234375,-0.0078125,0.03125,-0.0625,-0.0078125,-0.0234375,0.0234375,0.0078125,-0.0390625,0.0078125,0.015625,-0.0625,0.0234375,-0.0234375,0.2890625,-0.0625,-0.0234375,-0.0703125,0.0703125,-0.0234375,-0.03125,-0.15625,-0.0234375,0.0078125,-0.0078125,-0.0625,-0.015625,0.125,-0.140625,-0.1015625,0.0390625,0.0,0.109375,-0.0390625,-0.046875,-0.03125,0.0390625,0.078125,0.09375,-0.015625,0.0234375,0.0078125,-0.03125,0.140625,0.0859375,-0.03125,-0.1171875,-0.125,-0.0625,0.0390625,0.015625,0.1640625,0.0390625,-0.03125,-0.09375,0.015625,-0.03125,0.1171875,-0.0,-0.0625,0.0078125,-0.0078125,-0.078125,-0.0390625,0.0078125,-0.0390625,-0.0859375,-0.078125,0.0859375,-0.015625,0.0625,-0.0234375,-0.0390625,-0.03125,0.0625,-0.1328125,0.0234375,-0.015625,-0.0234375,0.0078125,-0.015625,-0.09375,0.046875,-0.1171875,-0.0546875,-0.0546875,0.125,0.2109375,0.1796875,-0.078125,-0.0078125,0.046875,-0.0859375,-0.0859375,-0.046875,-0.0,-0.0625,-0.015625,0.1015625,0.03125,-0.09375,-0.09375,-0.0234375,-0.1171875,-0.0390625,0.0625,-0.0703125,0.015625,-0.109375,-0.109375,-0.0234375,-0.0,0.0234375,0.1015625,0.078125,0.109375,-0.0,0.0703125,-0.0703125,0.171875,-0.03125,0.125,0.0078125,-0.046875,0.1015625,-0.0078125,-0.0703125,0.0234375,-0.0078125,-0.046875,0.0625,0.0546875,0.03125,-0.0234375,0.0078125,0.046875,0.0234375,-0.0078125,0.0859375,0.15625,-0.09375,-0.03125,0.046875,-0.03125,-0.0,-0.0078125,0.0,-0.0078125,0.0859375,0.0390625,-0.0234375,-0.0546875,-0.0859375,-0.0078125,0.0234375,-0.0390625,-0.015625,-0.0078125,0.1484375,-0.0390625,-0.0390625,0.0234375,-0.0,-0.0078125,0.0390625,-0.1171875,-0.0625,0.0546875,-0.03125,-0.0546875,-0.0234375,-0.0625,-0.0078125,0.0078125,-0.0,-0.0390625,0.0390625,0.015625,0.0,-0.03125,-0.0703125,0.015625,0.0078125,-0.0078125,0.0078125,-0.0234375,-0.03125,0.0,-0.0234375,-0.0078125,-0.0078125,-0.0,0.015625,-0.046875,0.0546875,-0.015625,0.0234375,0.046875,0.0,-0.1171875,-0.0390625,-0.03125,-0.0859375,-0.0234375,0.0234375,-0.03125,0.0234375,0.0546875,0.015625,0.0,-0.0859375,-0.0546875,0.0546875,0.0390625,0.03125,-0.0078125,-0.046875,-0.078125,0.1171875,0.0078125,0.0078125,-0.015625,0.015625,-0.015625,-0.015625,-0.0625,0.0234375,0.0,-0.0078125,0.0078125,0.0390625,0.0078125,-0.0390625,0.0078125,-0.015625,-0.0234375,0.0234375,0.125,0.015625,0.03125,0.0859375,0.0234375,-0.015625,-0.0234375,0.0078125,0.0234375,-0.0390625,0.0078125,-0.0625,-0.0078125,-0.1015625,-0.0234375,0.015625,-0.0078125,0.0625,-0.046875,-0.015625,-0.015625,-0.03125,0.03125,-0.015625,-0.0546875,-0.0234375,0.015625,-0.0390625,0.0625,-0.03125,0.015625,-0.0390625,0.0234375,-0.1328125,0.0390625,-0.0234375,-0.0625,0.015625,-0.1875,0.0390625,0.1171875,0.203125,-0.03125,0.046875,-0.1953125,0.0078125,-0.140625,0.0859375,-0.0703125,0.0546875,0.2265625,0.171875,0.0703125,-0.0234375,-0.234375,0.0390625,-0.015625,0.0390625,-0.0078125,0.0078125,0.0078125,0.0703125,0.015625,0.0078125,-0.15625,0.03125,0.0078125,0.046875,-0.015625,0.0546875,-0.1640625,0.1640625,-0.03125,-0.125,0.3046875,-0.015625,-0.0625,0.0390625,-0.0625,-0.1640625,-0.09375,0.078125,0.0,0.09375,0.0859375,-0.1015625,-0.0859375,-0.046875,0.0546875,-0.015625,-0.03125,-0.09375,-0.1796875,-0.078125,0.0,0.0078125,-0.09375,0.109375,0.0546875,-0.15625,0.140625,-0.0625,-0.03125,0.0234375,-0.078125,0.015625,-0.046875,0.1328125,0.09375,0.0,-0.1484375,0.078125,-0.09375,-0.09375,-0.0625,-0.1015625,0.0703125,-0.0625,-0.1328125,-0.109375,-0.015625,0.09375,-0.078125,-0.0078125,0.078125,-0.0859375,-0.1171875,0.0546875,0.1171875,-0.03125,0.0234375,0.0625,0.0390625,0.1171875,-0.046875,0.0078125,0.0078125,-0.1171875,-0.0234375,0.0234375,0.0546875,-0.0859375,0.03125,0.0859375,0.09375,-0.1171875,0.0703125,0.2109375,0.1875,0.015625,0.0,-0.0,-0.0078125,-0.1328125,-0.140625,-0.140625,0.046875,0.109375,0.1015625,-0.0625,-0.0234375,-0.0078125,-0.015625,0.0078125,-0.0,0.0078125,-0.0078125,-0.0,-0.0078125,-0.0078125,0.015625,0.0078125,-0.0,-0.0234375,-0.0234375,0.015625,-0.015625,-0.015625,-0.0078125,-0.0,0.0,-0.015625,-0.015625,0.015625,0.0,-0.015625,0.0,0.0,0.0078125,-0.0078125,0.0078125,-0.0078125,-0.0078125,-0.015625,-0.0,0.0078125,-0.0,-0.0,-0.0078125,-0.015625,0.015625,-0.015625,-0.0078125,-0.0078125,-0.0,0.0078125,-0.0078125,0.0,0.0078125,-0.0078125,0.0,-0.015625,-0.0,-0.0078125,-0.0078125,0.0,0.0,-0.0078125,0.0078125,0.0078125,-0.015625,-0.015625,0.0,-0.0,-0.0078125,-0.0078125,-0.0078125,0.0078125,-0.015625,0.015625,0.0078125,-0.0078125,-0.015625,-0.015625,-0.0078125,0.0,-0.0078125,-0.015625,-0.0078125,0.0,0.0,-0.0,-0.015625,-0.015625,-0.0234375,-0.0078125,-0.0,0.0,-0.015625,-0.015625,0.0078125,-0.0078125,0.0078125,-0.0,-0.0078125,-0.0078125,-0.0234375,-0.015625,0.0,-0.0078125,0.015625,0.0,-0.0078125,0.0,-0.0078125,-0.0078125,-0.0078125,-0.0,-0.0078125,-0.0078125,0.0,0.0078125,-0.0,-0.0078125,-0.0,-0.0078125,0.0078125,0.0,0.0078125,-0.0078125,-0.0,-0.015625,-0.0,-0.015625,-0.0078125,0.0,-0.015625,-0.015625,-0.015625,0.0078125,0.0078125,-0.015625,-0.015625,0.0078125,-0.015625,-0.0234375,0.0078125,0.0,0.0078125,-0.0,0.0,0.015625,-0.0078125,-0.0,-0.0078125,-0.015625,-0.0,-0.0078125,-0.0078125,-0.015625,-0.015625,0.0078125,0.0,-0.0078125,0.015625,-0.0078125,-0.0,-0.0234375,-0.0,-0.015625,0.015625,0.0078125,0.0078125,-0.0078125,0.0078125,0.0,0.0078125,0.0234375,0.0078125,0.0,-0.015625,-0.0234375,0.0234375,-0.0,0.015625,0.0078125,0.015625,0.0078125,0.0,-0.0078125,-0.0,-0.0078125,-0.0078125,-0.0234375,0.0,0.0078125,0.015625,0.0078125,0.0078125,-0.0,-0.0078125,-0.0078125,-0.0,0.0,0.0078125,-0.015625,0.0078125,0.0078125,0.0078125,-0.015625,-0.0078125,-0.015625,0.015625,-0.015625,-0.015625,0.0,-0.0078125,0.0078125,0.015625,-0.015625,0.0078125,0.0078125,-0.0078125,-0.015625,-0.015625,0.0234375,0.03125,0.015625,-0.015625,0.0234375,0.015625,-0.015625,-0.0078125,-0.0,-0.0078125,-0.0234375,-0.015625,0.0546875,-0.0078125,-0.0078125,0.015625,0.0,0.015625,-0.0078125,-0.015625,0.015625,-0.0078125,0.0078125,0.0,-0.0,-0.0078125,-0.0,0.03125,0.0078125,0.015625,0.03125,0.0078125,0.0,-0.0,-0.0078125,-0.0,0.03125,-0.0078125,-0.015625,-0.0078125,0.0078125,0.078125,0.1171875,0.046875,-0.0,-0.03125,0.0078125,-0.015625,0.078125,0.015625,0.046875,-0.09375,-0.09375,-0.046875,-0.0625,0.0703125,-0.0,-0.0,0.078125,-0.046875,-0.0390625,0.0078125,-0.0703125,-0.0546875,-0.015625,0.0078125,0.015625,0.046875,0.015625,0.0625,0.0078125,0.0078125,-0.03125,-0.0078125,-0.0078125,0.0078125,0.078125,0.109375,-0.0546875,0.03125,-0.0546875,0.140625,-0.0078125,0.015625,0.125,0.1328125,-0.0390625,0.015625,-0.015625,-0.0390625,0.0859375,-0.0234375,0.0234375,0.0546875,0.0625,0.046875,0.015625,0.0546875,-0.03125,0.0390625,-0.0703125,0.046875,0.046875,-0.0078125,0.015625,-0.0703125,0.0,-0.046875,0.0,0.15625,-0.0078125,-0.0078125,0.0078125,-0.015625,0.1015625,0.046875,-0.078125,-0.0703125,-0.0078125,0.0078125,-0.03125,0.0078125,0.03125,-0.015625,-0.0078125,-0.03125,-0.0546875,-0.0078125,0.0078125,0.015625,-0.046875,-0.015625,0.0078125,-0.046875,0.015625,0.09375,-0.03125,-0.0078125,-0.0390625,0.046875,0.015625,-0.046875,-0.0390625,-0.015625,0.125,0.0390625,0.0234375,0.0625,-0.0625,0.0,-0.046875,-0.03125,-0.0390625,0.03125,0.15625,0.0390625,0.0234375,0.015625,0.0390625,-0.0390625,0.0,-0.0234375,0.046875,-0.0,-0.125,0.1328125,0.03125,-0.03125,-0.0390625,0.09375,0.0859375,0.1875,-0.046875,0.015625,-0.0234375,0.0703125,-0.1328125,-0.0234375,0.0234375,-0.15625,-0.171875,0.0078125,-0.0234375,-0.1015625,-0.078125,-0.0234375,-0.0703125,0.0,0.0546875,0.0703125,-0.03125,0.078125,-0.0390625,0.0078125,0.0390625,0.0,0.03125,0.03125,-0.09375,0.0859375,0.1875,-0.1015625,0.0390625,-0.1328125,-0.0390625,0.046875,-0.0625,0.2109375,-0.140625,0.09375,-0.0078125,-0.03125,-0.03125,-0.0546875,0.03125,-0.015625,-0.046875,-0.0625,-0.0625,-0.0390625,0.078125,-0.0078125,-0.171875,0.0625,0.171875,-0.1171875,-0.03125,-0.0546875,0.0078125,-0.0390625,-0.015625,-0.1171875,-0.0,0.0546875,-0.015625,0.1328125,-0.0390625,-0.0703125,0.0859375,0.09375,0.0234375,-0.015625,0.109375,-0.0859375,0.0390625,-0.046875,-0.0,-0.078125,0.140625,-0.0859375,-0.1015625,-0.0390625,0.015625,-0.140625,0.1015625,-0.015625,-0.09375,0.015625,-0.0703125,0.0390625,0.0078125,-0.0546875,-0.015625,-0.0546875,0.1875,0.0234375,0.1015625,-0.15625,0.0625,0.0234375,-0.1484375,-0.09375,-0.09375,0.15625,-0.140625,-0.109375,0.09375,0.0234375,-0.0859375,-0.1015625,-0.078125,-0.1953125,-0.0703125,0.0234375,0.0234375,-0.03125,-0.1171875,0.0390625,0.171875,-0.0703125,-0.0546875,-0.0703125,-0.078125,0.03125,-0.015625,-0.1015625,0.078125,0.0546875,0.015625,0.078125,-0.015625,-0.0234375,0.0078125,-0.0625,0.0546875,0.015625,-0.078125,-0.078125,0.0546875,-0.046875,0.0625,0.0,0.0546875,0.0078125,0.078125,0.0078125,-0.0234375,-0.0234375,-0.0078125,-0.0078125,0.109375,-0.0078125,-0.046875,-0.015625,0.0,-0.0234375,0.03125,0.1015625,-0.0,0.015625,0.09375,0.015625,0.015625,-0.046875,-0.0546875,0.078125,0.03125,-0.015625,0.046875,-0.0390625,0.0,-0.015625,-0.09375,-0.015625,-0.0859375,-0.078125,-0.0234375,0.03125,-0.015625,-0.0546875,-0.0234375,-0.0078125,-0.0,0.0703125,0.03125,-0.0078125,0.015625,0.0390625,0.015625,0.0,-0.015625,-0.0625,0.0234375,0.0234375,0.0078125,-0.0078125,0.015625,0.0078125,-0.0703125,-0.0,-0.0234375,0.015625,-0.0390625,-0.1328125,-0.15625,0.046875,0.0859375,-0.1484375,-0.03125,0.0546875,0.0078125,-0.0546875,0.0078125,-0.0,-0.0078125,-0.03125,-0.0234375,0.015625,0.0625,0.03125,-0.0078125,-0.046875,0.03125,0.03125,-0.0546875,-0.0546875,0.1015625,-0.0859375,-0.0546875,0.0234375,0.0546875,-0.078125,0.0390625,0.0546875,-0.1328125,-0.0,0.046875,0.0078125,-0.0078125,0.0546875,-0.0859375,-0.0546875,-0.03125,-0.0625,-0.140625,-0.015625,-0.0078125,-0.0625,-0.0859375,-0.0,-0.0390625,-0.0859375,-0.0703125,-0.0390625,-0.1015625,-0.046875,-0.1171875,-0.0703125,0.125,0.1640625,0.03125,-0.1015625,0.203125,0.1015625,0.0625,0.1484375,-0.0859375,-0.046875,0.1875,0.015625,0.015625,0.0078125,-0.1640625,-0.0234375,-0.0625,0.046875,0.1328125,-0.1015625,0.0703125,0.1953125,0.015625,-0.0078125,0.1640625,-0.0625,0.0859375,0.1328125,-0.171875,0.09375,-0.0,0.0703125,0.0234375,-0.078125,0.0390625,0.1328125,-0.0078125,-0.109375,0.109375,0.046875,-0.1328125,0.0234375,-0.0390625,-0.09375,-0.078125,0.109375,0.1640625,-0.140625,0.109375,0.0859375,0.0546875,-0.1328125,-0.0546875,0.0625,0.03125,-0.015625,-0.0859375,-0.0859375,-0.0078125,-0.078125,0.03125,-0.0859375,0.046875,-0.078125,-0.0078125,0.0078125,0.078125,-0.0234375,0.140625,0.078125,-0.0703125,-0.0,-0.1171875,-0.171875,0.2578125,0.0703125,-0.0703125,-0.0390625,-0.046875,-0.0546875,0.03125,-0.1328125,0.015625,-0.203125,0.1328125,-0.03125,-0.0078125,-0.1953125,-0.1328125,0.03125,0.2421875,0.078125,-0.0703125,-0.109375,-0.0078125,-0.0546875,-0.140625,0.0390625,-0.140625,-0.0703125,-0.0546875,0.0390625,0.0,0.0625,-0.1171875,0.03125,0.203125,0.1171875,0.1640625,-0.109375,0.0625,-0.0234375,0.125,-0.0625,0.0078125,-0.1015625,0.03125,0.125,-0.0625,-0.0234375,0.15625,0.078125,-0.0,-0.0078125,0.0390625,-0.0546875,-0.0390625,0.0234375,0.0,-0.0,-0.0,-0.0390625,0.046875,-0.015625,-0.0390625,0.0390625,0.046875,0.0078125,0.140625,0.0234375,0.0078125,-0.0078125,0.0859375,0.09375,-0.0078125,-0.0625,0.0390625,0.0234375,-0.0234375,0.03125,-0.0390625,0.0078125,0.0625,0.1015625,0.0078125,-0.046875,0.0234375,0.0078125,-0.015625,-0.03125,0.0546875,-0.015625,-0.015625,0.015625,0.1171875,0.015625,-0.015625,-0.0078125,0.1171875,-0.046875,-0.109375,0.03125,0.0078125,0.015625,0.0546875,0.09375,-0.0546875,0.0546875,0.0703125,0.0390625,0.03125,0.0234375,0.0625,0.0390625,0.0546875,-0.03125,-0.0390625,0.0,-0.0,-0.046875,-0.078125,-0.0,-0.0078125,-0.0078125,0.0,-0.015625,-0.0078125,0.1171875,-0.015625,0.0078125,0.03125,-0.0390625,0.015625,0.03125,-0.015625,-0.0234375,0.0,0.015625,-0.015625,-0.015625,-0.109375,0.0078125,0.078125,0.0078125,0.0703125,-0.0546875,-0.0390625,-0.0078125,-0.015625,0.03125,0.1015625,0.0,-0.015625,-0.0390625,-0.015625,-0.1484375,-0.0234375,0.0390625,-0.0703125,-0.0078125,0.015625,0.03125,0.0078125,-0.0078125,0.0,-0.015625,0.0078125,-0.03125,-0.0625,0.0078125,-0.0,0.1328125,-0.0078125,0.078125,0.015625,0.015625,-0.0234375,-0.0078125,-0.0703125,-0.0,-0.015625,-0.0546875,-0.1171875,-0.078125,0.0625,0.234375,0.046875,-0.0234375,-0.09375,-0.1796875,0.0234375,0.0390625,0.09375,0.0546875,-0.078125,-0.1171875,0.0546875,-0.078125,-0.015625,-0.109375,-0.0078125,0.0234375,-0.078125,-0.03125,0.1484375,0.09375,-0.2109375,-0.0703125,-0.0,-0.1015625,0.0078125,0.0703125,-0.0546875,0.140625,-0.0390625,0.0,0.1328125,0.1796875,-0.03125,0.046875,-0.09375,0.0078125,0.078125,-0.0546875,-0.1015625,0.0,-0.203125,0.1171875,0.125,0.0625,-0.1015625,-0.140625,0.0703125,0.0234375,0.1015625,0.109375,0.0234375,-0.1328125,-0.046875,0.1484375,0.03125,0.0546875,-0.015625,0.046875,0.0546875,0.046875,0.171875,-0.1171875,-0.0859375,-0.0234375,-0.0625,0.125,-0.140625,-0.1953125,-0.0078125,-0.0625,0.0234375,0.09375,-0.0078125,0.0234375,-0.109375,-0.09375,-0.1015625,-0.2890625,-0.0625,-0.03125,0.03125,-0.1484375,0.078125,-0.171875,-0.015625,0.1328125,0.09375,-0.15625,-0.046875,0.09375,0.03125,-0.09375,-0.015625,0.1328125,0.2265625,0.1640625,0.03125,0.078125,0.0390625,0.046875,0.0546875,-0.015625,-0.109375,0.140625,-0.2265625,-0.0625,-0.1796875,0.1953125,0.0546875,0.046875,-0.109375,-0.1640625,0.0234375,0.0390625,-0.140625,0.1796875,0.015625,-0.109375,0.0234375,-0.03125,-0.1328125,-0.0546875,-0.1171875,0.046875,-0.0703125,0.0078125,-0.03125,-0.0234375,-0.03125,0.046875,0.015625,0.015625,-0.0390625,-0.0234375,-0.0625,0.0390625,0.03125,0.0546875,-0.046875,-0.015625,-0.015625,0.0078125,-0.0625,0.0078125,0.0390625,0.0703125,0.09375,0.1796875,-0.0625,-0.0390625,-0.0078125,0.046875,0.0,0.0234375,0.0234375,-0.078125,0.046875,-0.015625,-0.0,-0.0,0.015625,0.015625,0.1171875,-0.03125,-0.1015625,-0.0546875,0.0546875,-0.109375,0.015625,-0.0390625,0.0390625,-0.0703125,-0.0390625,-0.0234375,0.0625,-0.03125,0.015625,-0.0078125,0.015625,0.0,-0.0078125,-0.0078125,-0.03125,-0.0234375,0.03125,-0.03125,0.0,0.0078125,0.03125,-0.03125,0.1015625,-0.0078125,-0.0234375,0.015625,0.0546875,-0.015625,-0.0546875,0.015625,0.0390625,0.0078125,-0.0234375,-0.0390625,-0.0234375,0.0078125,-0.0390625,-0.0078125,0.0234375,0.125,-0.03125,0.03125,0.015625,0.0,0.1015625,0.0078125,0.078125,-0.0625,-0.03125,0.0234375,-0.0,0.0390625,0.109375,0.0,0.125,-0.015625,-0.1171875,0.078125,0.0078125,-0.0,0.03125,0.0625,-0.0625,0.015625,0.015625,0.0,0.0234375,0.0078125,0.046875,0.0546875,-0.0859375,0.0390625,0.078125,-0.0390625,0.03125,0.0390625,0.015625,0.015625,-0.0078125,0.0078125,0.0390625,0.0234375,-0.03125,0.015625,-0.0234375,0.1171875,0.0703125,-0.015625,0.015625,0.1015625,0.015625,0.0078125,-0.0078125,-0.0703125,-0.0078125,-0.03125,-0.0078125,0.0234375,0.109375,0.078125,0.0234375,0.015625,-0.015625,-0.1171875,0.015625,-0.0703125,0.078125,0.125,-0.03125,-0.0546875,0.046875,0.0703125,0.0859375,-0.015625,0.0390625,-0.0546875,-0.0390625,0.1015625,0.015625,-0.015625,0.0703125,0.0546875,-0.0,0.03125,-0.015625,-0.046875,0.0,0.015625,-0.0234375,0.0234375,-0.0234375,0.09375,-0.0,-0.0859375,-0.046875,-0.0390625,-0.0703125,-0.0078125,0.109375,0.046875,-0.0546875,0.0390625,-0.03125,0.078125,-0.0078125,0.0078125,0.0,-0.0703125,-0.046875,-0.09375,0.0078125,-0.09375,-0.0234375,-0.015625,-0.078125,0.015625,0.03125,0.03125,0.1015625,-0.0390625,-0.0859375,-0.1328125,0.046875,0.03125,-0.015625,0.0625,0.078125,0.03125,-0.0390625,-0.0625,-0.0234375,-0.0390625,0.078125,0.03125,0.109375,0.09375,-0.0234375,-0.0390625,0.0390625,0.1328125,0.109375,-0.046875,-0.03125,-0.1171875,-0.0390625,-0.015625,-0.015625,-0.0546875,-0.015625,0.0078125,0.015625,-0.109375,-0.0390625,-0.03125,-0.0390625,-0.0234375,-0.0078125,-0.03125,-0.0703125,0.0234375,0.03125,-0.09375,0.03125,0.0859375,-0.078125,0.1484375,0.1015625,-0.09375,0.0390625,-0.0390625,-0.046875,0.03125,-0.0234375,-0.0078125,-0.03125,0.0234375,-0.015625,-0.0625,-0.0,-0.0703125,0.0703125,0.015625,0.0859375,-0.0234375,-0.03125,-0.0390625,-0.015625,0.015625,-0.015625,-0.0078125,0.046875,-0.03125,-0.015625,-0.046875,0.015625,-0.09375,0.0234375,-0.0234375,0.03125,-0.046875,-0.0078125,0.0546875,-0.0234375,-0.0078125,-0.0234375,0.0078125,0.0625,0.0546875,0.03125,-0.0859375,-0.0703125,0.0859375,0.0234375,0.09375,-0.015625,0.0,0.09375,-0.0,-0.0625,-0.015625,0.03125,-0.0234375,0.0703125,0.15625,-0.03125,0.1484375,0.0078125,0.0078125,0.046875,-0.0078125,-0.0,-0.0546875,-0.0859375,0.1640625,-0.046875,0.0234375,0.046875,-0.1875,-0.0234375,0.0859375,-0.015625,-0.0234375,0.0078125,0.0234375,-0.0546875,-0.0234375,0.0625,-0.0078125,-0.0390625,0.0078125,0.015625,-0.0078125,-0.0,0.03125,0.0078125,-0.0703125,0.0,-0.0390625,0.015625,0.0,-0.0703125,-0.046875,-0.03125,0.0546875,-0.015625,-0.0078125,0.0078125,0.1171875,0.0078125,0.015625,-0.09375,0.015625,-0.03125,-0.203125,-0.046875,0.09375,-0.0625,0.0703125,0.1015625,-0.0078125,0.1015625,-0.0078125,0.0703125,0.015625,-0.0,0.1171875,0.015625,0.015625,-0.078125,0.15625,-0.0234375,-0.0234375,-0.015625,0.0703125,0.0234375,-0.0,0.015625,-0.1015625,0.0234375,0.0234375,-0.1171875,-0.015625,0.03125,0.0234375,-0.109375,-0.0625,-0.0546875,-0.078125,-0.0078125,0.1796875,-0.0546875,0.09375,0.0,-0.0234375,0.078125,-0.1171875,-0.0,0.046875,0.03125,0.046875,-0.03125,0.140625,0.0703125,-0.0703125,-0.1484375,-0.1015625,-0.0078125,0.0,-0.015625,-0.0625,-0.015625,-0.1015625,-0.1328125,-0.0390625,0.0546875,-0.0703125,-0.0625,0.015625,0.09375,-0.0859375,-0.0703125,-0.0859375,0.1328125,0.140625,-0.0078125,0.0546875,0.0546875,0.125,-0.0078125,-0.09375,0.0234375,0.046875,0.046875,-0.0625,-0.109375,0.0078125,-0.0859375,0.0078125,-0.0625,0.03125,0.1015625,-0.1796875,0.1640625,-0.171875,-0.0625,0.0859375,0.0859375,0.1484375,0.046875,-0.0859375,0.046875,-0.0546875,-0.1015625,-0.03125,-0.0703125,0.0078125,0.1171875,-0.0390625,-0.046875,-0.078125,0.2421875,0.015625,0.046875,-0.0,0.1015625,0.1171875,0.0,-0.0078125,0.0234375,-0.0390625,0.0,0.0703125,-0.015625,0.0078125,-0.03125,-0.078125,0.109375,-0.09375,0.0,-0.046875,-0.03125,-0.0078125,-0.1328125,-0.0859375,-0.0390625,0.015625,-0.015625,0.015625,0.0703125,-0.1484375,0.0234375,0.078125,-0.0703125,0.03125,-0.1484375,-0.0078125,0.1015625,-0.0546875,0.0546875,0.078125,-0.109375,-0.0,0.0078125,0.046875,0.0546875,-0.078125,-0.0,-0.0078125,0.0546875,0.015625,-0.0234375,0.03125,0.0078125,-0.015625,0.0,-0.0234375,-0.015625,0.03125,0.15625,-0.03125,-0.046875,0.0234375,-0.0234375,0.0234375,0.0078125,0.0,0.0234375,-0.0234375,0.0390625,-0.046875,-0.109375,-0.015625,0.0390625,0.09375,-0.0234375,-0.03125,0.0078125,0.015625,-0.015625,0.0859375,0.03125,0.0078125,-0.03125,0.0078125,-0.0,0.0546875,-0.0078125,0.078125,-0.03125,0.203125,0.0234375,0.1015625,0.0078125,-0.0078125,0.0546875,-0.015625,0.0,-0.0,-0.0234375,-0.0390625,-0.078125,-0.0078125,-0.078125,0.0859375,0.0,-0.015625,0.0078125,-0.0703125,0.0234375,0.015625,-0.0234375,-0.015625,-0.0078125,-0.0,-0.0078125,-0.0390625,0.0078125,-0.015625,0.015625,-0.078125,-0.046875,-0.09375,-0.015625,-0.015625,-0.0390625,-0.03125,-0.046875,0.046875,0.0078125,-0.0859375,0.0,-0.0859375,0.0546875,-0.0390625,0.015625,0.0078125,-0.03125,-0.0859375,-0.109375,-0.0078125,0.0078125,0.0078125,-0.0078125,-0.03125,0.0234375,-0.0078125,0.0078125,-0.015625,0.09375,-0.03125,-0.015625,-0.0078125,-0.0546875,0.0,-0.0078125,0.0625,-0.109375,-0.0078125,0.078125,-0.0078125,-0.0234375,-0.015625,0.15625,0.09375,0.1328125,-0.0234375,-0.0546875,-0.0390625,0.0,0.0234375,-0.0390625,-0.015625,-0.015625,-0.046875,0.046875,0.0390625,-0.0859375,0.0,0.03125,-0.078125,0.046875,-0.0234375,-0.03125,0.0625,0.046875,0.1171875,0.0078125,0.0546875,-0.0625,-0.03125,0.0703125,-0.0,0.078125,-0.078125,0.0,0.0390625,0.03125,-0.0703125,0.015625,-0.0546875,-0.015625,-0.0390625,-0.03125,0.078125,0.03125,-0.0546875,0.0234375,0.0625,-0.046875,-0.0234375,-0.0703125,0.1015625,0.0078125,0.046875,0.0,-0.0390625,-0.0,-0.0078125,-0.0390625,-0.0390625,0.0,0.03125,0.078125,-0.0234375,0.03125,0.125,0.0078125,0.0078125,0.046875,-0.0234375,-0.046875,0.0234375,-0.0703125,0.0,0.015625,-0.0078125,-0.09375,-0.09375,0.03125,0.125,-0.015625,0.0546875,-0.0546875,0.0,-0.0703125,0.015625,0.046875,0.0078125,-0.03125,0.0078125,-0.0703125,-0.0625,-0.0234375,0.046875,-0.0546875,-0.0390625,0.0390625,-0.046875,-0.078125,0.0390625,-0.0078125,-0.0,-0.0078125,0.0,0.0078125,0.015625,0.0625,-0.09375,0.046875,0.0390625,-0.0546875,-0.0,-0.015625,-0.0078125,0.0078125,-0.078125,0.0703125,0.03125,-0.0546875,-0.0859375,0.0703125,-0.15625,-0.0546875,0.1015625,0.0,-0.03125,-0.1015625,-0.046875,0.0234375,-0.03125,0.0390625,0.046875,0.0078125,-0.0859375,-0.03125,-0.0625,-0.0078125,-0.0390625,0.0234375,-0.0078125,-0.0078125,-0.046875,-0.0390625,-0.03125,-0.0078125,-0.015625,0.0234375,0.015625,0.0,0.0,0.015625,-0.015625,0.0078125,0.0390625,-0.0546875,0.0,-0.0,-0.0390625,0.0859375,0.015625,0.0,0.0078125,0.0234375,-0.0390625,-0.015625,-0.0234375,-0.0078125,-0.0234375,-0.0078125,-0.0078125,0.0,0.03125,-0.015625,-0.015625,0.015625,-0.0390625,0.0,0.0078125,-0.015625,-0.015625,0.03125,0.0859375,-0.0703125,0.0390625,0.09375,0.0390625,0.03125,0.0859375,-0.0390625,0.09375,-0.015625,0.03125,0.0390625,-0.0234375,0.03125,0.0078125,0.0390625,-0.015625,-0.0234375,0.015625,-0.0078125,0.0546875,-0.0078125,0.015625,-0.03125,0.0546875,0.0234375,-0.0078125,-0.0078125,0.046875,0.0078125,-0.0390625,-0.0,0.03125,-0.0234375,0.0234375,-0.0,0.0,-0.0234375,0.015625,0.0078125,-0.015625,-0.0078125,0.015625,0.0703125,-0.1328125,0.015625,-0.0546875,-0.015625,-0.0546875,0.0390625,0.0,-0.015625,0.015625,-0.0390625,0.015625,0.015625,0.015625,-0.0078125,-0.0,-0.0234375,0.078125,-0.0,0.0859375,0.0546875,-0.03125,-0.0078125,-0.0234375,0.0703125,-0.0390625,-0.0546875,-0.0078125,-0.0625,-0.0078125,-0.0234375,-0.0078125,0.015625,-0.0234375,0.0,-0.0703125,0.015625,-0.03125,-0.109375,0.0234375,0.0078125,-0.015625,0.0,-0.0,0.0,0.0859375,0.0078125,-0.046875,-0.0234375,-0.03125,-0.0625,0.09375,0.0703125,-0.0078125,-0.046875,-0.0390625,-0.0234375,0.046875,-0.0078125,-0.0,0.015625,-0.0625,-0.078125,-0.03125,-0.046875,-0.0078125,0.015625,0.0234375,-0.0,-0.0,-0.046875,-0.0,0.046875,0.0234375,-0.0625,0.0078125,-0.0390625,-0.109375,-0.0546875,0.0,-0.0703125,0.0625,0.0703125,0.0390625,-0.0390625,-0.0625,0.03125,0.0234375,0.0625,0.0,0.03125,-0.0234375,0.0,0.0,-0.0390625,-0.015625,0.0546875,0.03125,0.140625,0.0078125,0.0,0.015625,0.0390625,-0.046875,-0.078125,0.03125,0.0234375,0.046875,0.0234375,-0.015625,0.0,0.0546875,-0.0546875,-0.0390625,-0.0703125,0.015625,-0.0,0.0078125,0.0234375,-0.0078125,0.109375,-0.0078125,-0.0,-0.0859375,-0.0546875,-0.03125,0.0703125,-0.0234375,-0.046875,0.0,0.015625,0.015625,-0.0390625,0.015625,-0.0078125,-0.0546875,-0.0234375,-0.0234375,0.0234375,0.0234375,0.03125,-0.015625,0.0078125,0.03125,-0.03125,0.015625,-0.015625,0.015625,0.0546875,-0.0,-0.046875,-0.046875,-0.0703125,0.109375,-0.0078125,0.0234375,-0.0703125,-0.03125,0.046875,-0.0625,-0.0390625,0.0390625,0.0546875,-0.0625,-0.046875,0.0390625,-0.0625,-0.0078125,-0.0078125,-0.0,0.0546875,0.0546875,-0.015625,0.1015625,-0.0390625,-0.03125,-0.0078125,0.078125,-0.015625,-0.0,0.03125,-0.0546875,0.0078125,-0.015625,-0.0078125,0.0,0.0234375,-0.0390625,-0.0,-0.03125,-0.0703125,0.1015625,0.015625,-0.0078125,-0.03125,0.015625,-0.0078125,-0.078125,0.03125,-0.03125,-0.0078125,-0.0,0.03125,-0.0,0.0,0.0078125,-0.03125,0.046875,-0.0078125,-0.015625,0.0234375,-0.0,0.0078125,0.0703125,-0.09375,0.015625,-0.0390625,0.0625,0.078125,0.03125,0.015625,-0.015625,0.0078125,0.03125,0.0078125,0.0390625,0.0859375,-0.03125,0.0234375,-0.0078125,-0.03125,0.0078125,-0.0234375,-0.046875,0.03125,0.0234375,-0.046875,0.015625,0.015625,0.0234375,-0.0546875,0.03125,-0.015625,-0.0390625,-0.0078125,0.125,-0.0546875,0.0,-0.078125,-0.03125,-0.0234375,0.0078125,-0.03125,-0.0390625,0.0078125,0.015625,0.0078125,-0.0234375,0.0078125,-0.078125,0.03125,0.09375,0.015625,0.0078125,-0.0,0.015625,0.046875,-0.015625,0.0078125,-0.015625,-0.015625,-0.015625,0.0078125,-0.0078125,-0.0703125,-0.0078125,0.015625,-0.0078125,-0.0234375,-0.0703125,0.0546875,0.015625,0.0,-0.015625,0.0078125,-0.0078125,-0.03125,-0.0234375,-0.03125,-0.046875,0.0234375,0.0390625,0.0078125,-0.0078125,-0.015625,-0.0546875,0.0078125,0.0234375,0.0625,0.015625,-0.0234375,-0.0546875,0.0390625,-0.0,-0.0234375,-0.0078125,0.0703125,0.046875,-0.0234375,-0.0234375,-0.0390625,-0.1328125,0.0625,-0.0078125,0.0390625,0.0078125,-0.046875,-0.0390625,0.015625,0.171875,-0.03125,-0.0703125,0.0234375,-0.0703125,-0.078125,0.046875,0.0078125,0.0546875,0.015625,0.09375,0.21875,-0.109375,-0.078125,-0.0703125,-0.0703125,-0.046875,-0.0234375,0.0078125,-0.0078125,-0.0078125,0.046875,0.0625,-0.0625,0.0234375,-0.0703125,0.09375,-0.015625,-0.0234375,-0.046875,-0.1015625,-0.0625,0.1171875,-0.0390625,0.0,0.046875,-0.0625,0.0078125,0.078125,0.0234375,-0.09375,-0.09375,-0.03125,0.15625,-0.046875,0.046875,0.140625,0.03125,-0.0078125,0.0625,-0.046875,-0.0859375,-0.0078125,0.0625,0.046875,-0.046875,0.0234375,0.0078125,0.0234375,-0.015625,-0.0,-0.0390625,0.21875,-0.0234375,0.0390625,-0.015625,-0.0625,-0.0,-0.0234375,0.03125,-0.0234375,0.0390625,-0.0546875,-0.0234375,0.0859375,-0.09375,0.0546875,-0.046875,0.015625,-0.0078125,-0.109375,-0.0546875,0.0859375,0.0703125,0.203125,-0.0078125,-0.046875,0.1328125,0.125,0.0234375,-0.0546875,-0.0390625,-0.0859375,-0.0234375,0.15625,0.015625,-0.046875,0.0234375,-0.03125,0.0078125,-0.21875,-0.0234375,-0.046875,-0.0,0.125,-0.03125,0.015625,-0.1484375,0.046875,-0.078125,-0.0078125,-0.03125,-0.0390625,-0.0078125,-0.0234375,0.0390625,0.0234375,-0.015625,-0.0234375,-0.0078125,-0.03125,0.1015625,-0.0234375,-0.0078125,-0.0078125,0.0546875,-0.09375,-0.1015625,-0.03125,-0.0234375,0.0,0.046875,0.125,0.0234375,-0.0859375,0.0546875,-0.0,0.0078125,-0.0546875,-0.0234375,-0.03125,-0.09375,-0.0078125,-0.0234375,0.03125,0.046875,-0.0078125,0.0703125,0.046875,0.0859375,-0.0859375,0.015625,-0.0390625,-0.0859375,-0.0546875,-0.0,-0.0625,0.0703125,-0.0234375,-0.15625,-0.03125,-0.03125,0.015625,-0.0703125,-0.0234375,-0.015625,0.0,0.09375,-0.015625,0.046875,0.046875,0.015625,-0.03125,-0.0,-0.015625,-0.0078125,-0.03125,0.078125,-0.1171875,-0.03125,0.0859375,-0.0390625,-0.015625,0.140625,0.0390625,0.0078125,0.1015625,0.0078125,0.0078125,-0.0,-0.0234375,-0.015625,0.015625,-0.0,0.03125,0.0,-0.03125,-0.03125,-0.0390625,-0.046875,0.015625,-0.03125,-0.078125,0.09375,-0.0,-0.0078125,-0.0078125,0.0078125,0.0625,0.0390625,-0.0234375,-0.015625,-0.0625,-0.0859375,-0.1015625,-0.0390625,-0.078125,-0.0078125,-0.078125,0.078125,-0.046875,0.03125,0.0,0.125,0.046875,-0.0390625,-0.03125,0.0234375,-0.03125,-0.03125,0.0703125,-0.0078125,-0.0390625,-0.015625,0.0078125,0.0078125,-0.0,-0.046875,0.0078125,-0.0078125,-0.0390625,-0.0703125,0.1875,0.0625,-0.03125,-0.125,0.09375,-0.15625,0.0390625,-0.0078125,0.0234375,0.1328125,-0.078125,0.0625,0.0703125,-0.0234375,0.0625,-0.0859375,0.0234375,0.234375,-0.0078125,-0.0234375,-0.140625,0.0078125,0.0546875,-0.1171875,0.0390625,-0.0390625,0.015625,-0.015625,0.03125,0.1484375,-0.125,0.078125,-0.1171875,0.046875,0.015625,0.3046875,0.125,0.171875,0.1328125,-0.109375,-0.03125,-0.09375,0.015625,0.015625,0.015625,-0.0234375,0.046875,-0.015625,0.0703125,-0.09375,-0.0390625,0.140625,0.03125,0.09375,0.1796875,0.0546875,-0.0546875,-0.0703125,-0.078125,0.03125,0.0078125,-0.125,0.0234375,0.0,0.03125,0.046875,0.0390625,0.109375,0.0234375,-0.0390625,-0.140625,0.078125,-0.03125,-0.078125,0.09375,-0.0234375,0.0,0.0703125,0.0078125,0.140625,0.109375,-0.140625,-0.0,0.0234375,0.21875,-0.0,-0.046875,-0.078125,0.140625,-0.0859375,0.0546875,-0.0625,0.046875,-0.03125,-0.015625,0.0078125,-0.109375,0.0625,-0.015625,-0.0859375,0.09375,-0.09375,0.09375,0.0234375,0.0,0.03125,0.2109375,0.1015625,-0.078125,0.0546875,-0.109375,0.0390625,-0.1328125,0.046875,-0.09375,0.0390625,0.0625,0.2109375,-0.0234375,0.0078125,0.125,-0.09375,0.125,0.125,0.0390625,0.0390625,-0.015625,-0.046875,-0.03125,0.015625,0.0546875,-0.0546875,0.0546875,0.0078125,-0.03125,0.0625,-0.015625,0.015625,-0.046875,0.0078125,0.0,-0.046875,-0.09375,-0.0078125,0.0078125,0.0390625,-0.0234375,-0.0078125,0.0234375,-0.0390625,0.0625,0.0390625,-0.046875,0.0078125,-0.046875,0.0234375,0.0078125,-0.0078125,-0.03125,-0.03125,0.03125,-0.0234375,0.0234375,0.0546875,-0.0625,0.0234375,0.015625,-0.0,-0.0859375,-0.0546875,-0.0390625,0.0546875,0.0546875,-0.015625,0.0078125,0.046875,0.015625,0.015625,-0.0546875,-0.015625,0.0078125,0.0390625,-0.0390625,0.0,0.0859375,-0.046875,-0.0234375,0.015625,0.0390625,-0.015625,-0.0,0.03125,0.0234375,-0.0234375,-0.0234375,-0.0078125,0.03125,0.0,-0.0625,0.0390625,0.0546875,0.0,-0.0,-0.0234375,0.0234375,0.0390625,0.0078125,-0.046875,-0.0859375,-0.0234375,-0.0625,-0.0390625,-0.015625,-0.0390625,0.0,-0.03125,-0.046875,0.0234375,-0.046875,0.0,0.0,-0.0078125,0.0078125,0.03125,0.0,-0.0078125,0.03125,-0.0078125,0.03125,-0.0625,-0.0234375,-0.03125,0.0078125,-0.109375,0.0,-0.0625,-0.03125,-0.0234375,0.03125,0.0078125,0.0390625,0.0234375,-0.0546875,-0.015625,0.0234375,-0.078125,0.0078125,0.0,-0.0234375,0.0234375,0.0078125,0.0,0.046875,-0.0,-0.03125,-0.0078125,0.03125,-0.0703125,-0.0703125,-0.171875,-0.109375,0.1328125,-0.015625,0.0234375,-0.0390625,0.0078125,0.0390625,0.1015625,-0.0390625,-0.109375,0.046875,0.3359375,-0.09375,0.140625,-0.0546875,-0.078125,0.0546875,-0.140625,0.0546875,0.0078125,0.1171875,-0.1015625,-0.046875,-0.078125,0.0078125,-0.0703125,0.0859375,0.125,0.03125,-0.078125,-0.078125,0.1171875,-0.0703125,0.0,-0.1484375,-0.1328125,0.015625,-0.0234375,0.1015625,0.171875,-0.0546875,-0.046875,0.03125,0.0703125,-0.1015625,0.125,0.09375,-0.0078125,0.0703125,-0.1015625,-0.0546875,-0.0703125,-0.140625,0.03125,0.0078125,0.140625,0.1640625,0.1640625,0.1171875,0.1328125,-0.0859375,0.03125,0.15625,0.0546875,0.03125,-0.0546875,-0.09375,0.046875,-0.0078125,0.015625,-0.0390625,-0.0390625,-0.1171875,-0.046875,-0.03125,0.0703125,-0.09375,-0.1015625,-0.03125,-0.0625,0.0859375,-0.09375,0.078125,-0.140625,0.15625,0.0703125,0.015625,0.0625,0.0703125,0.046875,-0.109375,0.109375,0.0234375,-0.1484375,0.0234375,-0.0078125,0.046875,-0.0859375,0.0,0.1171875,0.0078125,-0.015625,-0.140625,0.0078125,-0.1015625,0.15625,0.0625,-0.03125,-0.0078125,0.1171875,-0.0078125,-0.09375,0.0078125,-0.0546875,0.1015625,0.25,-0.0546875,0.1171875,0.0234375,-0.0625,0.0703125,-0.0625,0.1328125,0.1328125,-0.0234375,0.0,0.0,0.0,-0.0078125,-0.0078125,0.0078125,-0.0078125,-0.0078125,-0.0234375,-0.0234375,0.015625,-0.0234375,0.015625,-0.046875,-0.015625,-0.015625,0.03125,0.0,-0.03125,0.0078125,-0.03125,-0.03125,0.015625,-0.015625,-0.03125,0.0,-0.0078125,-0.015625,-0.0078125,-0.015625,0.0,-0.015625,0.0078125,-0.0,-0.0234375,-0.0234375,-0.0234375,-0.0234375,-0.0234375,-0.0390625,0.0078125,0.0234375,0.0,-0.0,0.015625,-0.0234375,-0.0,-0.015625,-0.0625,-0.015625,0.03125,0.0,-0.03125,0.0,0.0,0.0625,-0.0078125,-0.015625,-0.0,0.0,-0.0078125,-0.015625,-0.0234375,0.0234375,0.0,0.0234375,0.0078125,-0.0234375,-0.0390625,0.0,0.0078125,0.0234375,-0.015625,-0.0078125,-0.0078125,-0.0078125,-0.015625,-0.0,0.0234375,0.0,-0.0078125,-0.0,0.015625,-0.03125,-0.0078125,-0.015625,-0.0234375,0.0,-0.0390625,-0.015625,-0.0234375,0.015625,0.0,-0.0,-0.03125,-0.0390625,-0.0078125,0.015625,0.0078125,-0.046875,-0.015625,0.015625,0.0,-0.0234375,0.0546875,-0.0078125,0.0078125,-0.0,-0.015625,-0.0234375,-0.015625,0.0625,-0.03125,-0.0234375,-0.0234375,-0.0078125,-0.03125,-0.0078125,-0.015625,-0.0234375,-0.015625,0.0,0.0234375,-0.0234375,-0.015625,0.0078125,0.0390625,0.0078125,-0.0078125,0.015625,-0.0,0.0078125,-0.015625,-0.0078125,0.0078125,-0.0625,0.0390625,-0.0078125,0.0078125,-0.015625,0.0234375,0.0234375,0.03125,0.046875,0.0703125,0.015625,0.0078125,0.0,-0.0234375,-0.015625,0.0078125,0.015625,-0.0078125,-0.015625,0.03125,0.03125,-0.03125,0.0234375,0.0234375,-0.0234375,0.015625,-0.0234375,0.0,0.0078125,0.0234375,-0.0078125,-0.0390625,0.0546875,-0.015625,0.0078125,0.0546875,-0.0234375,-0.015625,0.0390625,-0.015625,0.03125,-0.03125,0.0078125,-0.0078125,0.046875,-0.0234375,-0.0234375,-0.046875,-0.0078125,-0.0,-0.0390625,-0.0234375,-0.0234375,-0.03125,0.015625,0.0390625,0.0234375,0.0234375,0.015625,0.0078125,0.0078125,-0.0078125,-0.0,-0.03125,0.0078125,-0.0234375,-0.0,-0.0078125,0.015625,0.0078125,0.015625,-0.046875,-0.0078125,-0.0078125,0.015625,-0.0234375,0.015625,-0.015625,0.0078125,-0.0078125,0.0,-0.0078125,-0.0078125,0.0390625,0.0078125,-0.0078125,-0.03125,0.0078125,-0.03125,-0.015625,-0.0234375,-0.0234375,-0.015625,0.0234375,0.015625,-0.03125,0.015625,-0.0078125,0.0234375,-0.0390625,-0.0078125,-0.0390625,-0.0078125,-0.0234375,0.015625,-0.0234375,-0.0,0.0078125,-0.03125,-0.0234375,-0.0078125,-0.0078125,0.0078125,0.0234375,0.0546875,0.0234375,0.0078125,0.078125,-0.0,0.0390625,-0.03125,0.0,0.015625,0.0,-0.0078125,-0.0,0.015625,-0.015625,-0.0234375,0.015625,-0.0078125,-0.015625,-0.015625,-0.0234375,0.0859375,-0.0234375,0.0,-0.0546875,-0.015625,0.0078125,0.0,-0.03125,0.0,0.015625,0.0625,-0.015625,0.015625,0.0,0.0078125,0.0078125,-0.0078125,0.03125,0.0,0.0234375,-0.015625,-0.0390625,0.0234375,0.0625,-0.046875,-0.0546875,0.0859375,0.0390625,0.0546875,0.03125,-0.0078125,0.0078125,-0.0,-0.0546875,-0.0234375,0.0234375,-0.0078125,0.0,0.0,-0.0078125,0.03125,-0.0078125,-0.0234375,-0.0078125,-0.015625,0.0390625,-0.0390625,0.0,0.0234375,-0.03125,-0.0,-0.0234375,-0.0234375,-0.015625,-0.0390625,-0.078125,0.0,0.0546875,-0.0234375,-0.0234375,0.015625,-0.0078125,-0.0234375,-0.0078125,0.0078125,0.0078125,0.0390625,-0.0078125,-0.015625,0.0234375,-0.0390625,0.0234375,-0.0078125,-0.0078125,0.0078125,-0.078125,-0.0,-0.0078125,-0.0,0.015625,-0.015625,-0.015625,-0.0703125,-0.015625,-0.0,-0.0390625,-0.03125,-0.0,-0.03125,-0.0234375,-0.0,-0.0234375,-0.015625,0.03125,0.0078125,-0.0234375,-0.0078125,-0.015625,-0.015625,0.09375,0.0703125,0.046875,0.0234375,0.0625,-0.0,0.0078125,-0.015625,-0.0234375,0.0078125,-0.0078125,0.0078125,0.03125,-0.0078125,0.03125,-0.0,0.1171875,-0.0078125,0.0703125,-0.046875,-0.0234375,-0.0703125,-0.0390625,-0.046875,-0.0859375,0.109375,-0.0234375,0.1171875,0.0546875,-0.015625,-0.1015625,-0.0,-0.1328125,0.0,0.015625,-0.078125,-0.0078125,-0.03125,0.1015625,-0.015625,0.0078125,0.015625,-0.0,0.0703125,-0.03125,-0.046875,-0.078125,0.0234375,-0.046875,0.0859375,-0.0703125,0.0,0.0546875,0.015625,0.0546875,-0.0,0.09375,-0.078125,-0.0078125,0.1953125,-0.0390625,-0.03125,0.125,0.015625,0.0546875,-0.03125,-0.0078125,-0.0390625,0.015625,0.0234375,0.1328125,-0.0078125,-0.0390625,0.015625,-0.0,-0.1015625,0.0078125,0.1015625,-0.078125,-0.015625,-0.078125,-0.1171875,-0.0390625,-0.09375,0.046875,0.2890625,-0.0390625,0.0078125,0.0625,-0.0390625,0.0,-0.0078125,0.0234375,0.015625,0.0,0.0390625,-0.03125,-0.0078125,-0.078125,-0.0390625,0.0546875,0.0234375,0.078125,-0.0625,0.0078125,-0.0546875,0.0390625,-0.0625,-0.03125,0.015625,-0.0390625,-0.0078125,-0.0625,0.0234375,0.046875,-0.0,0.0078125,0.015625,0.0546875,0.0703125,-0.046875,-0.046875,0.03125,0.0625,0.0234375,-0.015625,0.0703125,-0.015625,-0.015625,0.03125,0.0,0.09375,0.03125,-0.0,-0.0390625,-0.078125,0.015625,-0.0625,-0.0078125,-0.015625,0.03125,-0.046875,-0.015625,0.0390625,0.0390625,0.03125,0.015625,0.0234375,0.015625,0.03125,0.015625,-0.015625,0.0,0.046875,-0.0234375,0.0390625,-0.0234375,0.0625,0.046875,-0.0078125,0.015625,-0.0546875,0.0,0.0078125,-0.046875,-0.0625,0.0234375,-0.0546875,0.0703125,-0.0078125,0.125,-0.015625,-0.03125,0.1015625,0.0078125,0.0078125,0.0078125,0.0078125,-0.0234375,-0.046875,0.0078125,0.0078125,0.0,-0.015625,-0.0546875,0.0078125,-0.0625,0.109375,0.1015625,0.03125,0.0234375,-0.0078125,-0.03125,0.0390625,0.0,0.03125,-0.046875,-0.0078125,-0.046875,-0.03125,-0.03125,-0.046875,-0.0234375,0.0234375,0.0390625,0.0078125,-0.046875,0.0703125,-0.0546875,-0.0703125,0.0,0.0546875,-0.046875,-0.046875,0.0234375,-0.0390625,-0.0,-0.0078125,-0.0234375,0.0234375,0.0234375,-0.0234375,-0.015625,0.1484375,0.0078125,-0.0,-0.046875,0.0546875,0.0390625,-0.015625,-0.1328125,0.0078125,-0.09375,0.03125,0.1015625,-0.0078125,-0.015625,-0.0390625,-0.046875,-0.03125,-0.0625,-0.0078125,0.0859375,0.109375,0.0703125,-0.0703125,0.0078125,-0.03125,0.015625,-0.046875,0.0859375,-0.0078125,0.0,-0.015625,-0.015625,0.0234375,0.0546875,-0.0390625,-0.0234375,0.015625,-0.0234375,-0.0390625,-0.0078125,-0.0546875,0.0078125,0.0,-0.03125,-0.078125,-0.0234375,0.0234375,0.0,-0.0,-0.0234375,-0.0234375,0.046875,0.3046875,-0.03125,0.0625,-0.0234375,-0.078125,0.015625,-0.109375,0.1015625,-0.09375,-0.0234375,-0.0078125,-0.140625,0.0703125,0.09375,0.0625,0.0234375,0.0703125,0.171875,-0.046875,0.078125,-0.1171875,-0.0625,-0.1015625,-0.03125,-0.0546875,0.0234375,0.015625,-0.046875,-0.0859375,-0.078125,0.078125,0.046875,0.109375,-0.046875,0.1015625,0.046875,-0.109375,0.078125,-0.0078125,0.03125,0.0703125,-0.03125,-0.0078125,0.109375,0.109375,-0.1015625,-0.046875,-0.0390625,-0.03125,0.109375,0.1015625,-0.0390625,0.078125,0.2109375,-0.0234375,-0.046875,0.0234375,-0.0859375,-0.0078125,0.0234375,-0.1015625,0.0234375,-0.0546875,0.109375,0.015625,0.171875,-0.1171875,-0.0234375,-0.0,0.109375,0.109375,0.0234375,-0.078125,0.0546875,0.03125,-0.078125,0.0546875,0.109375,-0.0859375,-0.1171875,-0.015625,-0.109375,-0.015625,-0.15625,-0.1640625,-0.0859375,0.046875,0.09375,-0.078125,-0.015625,0.0625,-0.078125,0.0859375,0.0,-0.0078125,-0.046875,0.0703125,-0.0390625,-0.0078125,-0.03125,-0.0859375,0.0,0.03125,-0.0859375,0.0703125,-0.0546875,0.0078125,0.0546875,-0.0234375,0.0078125,0.0234375,0.0234375,-0.0625,0.0703125,0.0625,-0.109375,0.1640625,-0.0234375,-0.0390625,0.015625,0.0859375,0.0859375,0.03125,-0.046875,-0.0,-0.015625,0.1484375,-0.0078125,-0.0546875,-0.0078125,-0.015625,0.0234375,0.0078125,0.0390625,-0.015625,0.0,-0.078125,-0.0546875,0.0,0.0859375,0.0078125,0.0703125,0.0546875,0.0703125,-0.109375,-0.078125,0.0390625,-0.046875,0.0234375,0.078125,-0.046875,-0.015625,0.0078125,0.03125,-0.0078125,-0.03125,0.0078125,-0.0390625,0.1484375,0.09375,-0.015625,-0.0390625,0.1796875,-0.015625,0.03125,-0.0859375,-0.015625,0.0625,0.0546875,0.0390625,0.0234375,-0.0390625,-0.0234375,-0.0078125,0.0390625,-0.0703125,0.03125,-0.0546875,-0.015625,0.0078125,0.015625,-0.0078125,-0.0078125,-0.0,0.0390625,-0.0,-0.0234375,0.0625,-0.03125,-0.0,-0.1015625,-0.0078125,0.0546875,0.0859375,0.03125,-0.015625,0.015625,-0.0546875,-0.015625,-0.0390625,-0.1484375,-0.015625,0.0390625,-0.0234375,-0.0625,0.015625,-0.0078125,-0.0703125,0.0859375,-0.0,-0.0078125,0.03125,-0.0234375,0.0703125,-0.1015625,0.0546875,0.0234375,-0.0,0.1171875,0.046875,-0.0,0.015625,-0.0390625,0.046875,0.0234375,-0.0078125,0.0703125,0.0,-0.0,0.078125,-0.0078125,-0.0546875,0.015625,0.09375,-0.0,-0.0546875,-0.0234375,-0.0,0.0078125,0.0390625,0.140625,-0.0546875,-0.03125,-0.0078125,-0.0,0.09375,0.0078125,-0.109375,-0.0078125,0.09375,-0.046875,-0.0234375,0.046875,-0.0234375,-0.125,0.0703125,0.2421875,0.0078125,-0.109375,-0.0234375,-0.0625,0.09375,-0.09375,0.0703125,-0.078125,0.1171875,-0.0390625,-0.0859375,-0.0703125,-0.0546875,0.0,-0.1015625,0.015625,0.3359375,-0.0390625,0.0703125,0.0703125,0.171875,0.21875,-0.078125,0.03125,0.28125,-0.0546875,0.0625,-0.21875,-0.03125,0.0546875,-0.0234375,0.0546875,-0.078125,0.0234375,-0.0859375,-0.1328125,0.046875,0.125,-0.0625,-0.125,0.125,-0.0,-0.140625,-0.0234375,-0.0625,-0.171875,-0.046875,0.1640625,0.0859375,0.0,-0.046875,0.1015625,-0.0390625,-0.1171875,-0.0859375,-0.0234375,-0.0625,0.0859375,0.1015625,-0.0390625,0.09375,-0.1953125,0.25,0.203125,0.0546875,-0.0078125,0.1484375,0.0390625,-0.0390625,0.046875,-0.1015625,-0.0390625,0.0703125,-0.0078125,-0.109375,0.015625,-0.15625,-0.03125,-0.0078125,-0.0625,-0.1015625,0.015625,0.03125,0.1328125,-0.0625,-0.078125,-0.140625,0.0390625,0.0625,-0.015625,-0.0859375,-0.1796875,0.0390625,0.09375,0.0546875,-0.1328125,-0.078125,-0.234375,-0.0234375,-0.1484375,0.1640625,0.09375,0.0078125,0.0234375,-0.09375,-0.046875,-0.109375,-0.03125,0.0,0.0,0.046875,0.1484375,0.2265625,-0.0078125,0.0546875,0.2265625,-0.140625,-0.03125,-0.09375,0.0078125,-0.09375,0.09375,-0.03125,0.03125,0.0390625,0.03125,0.0546875,-0.0,-0.0,0.03125,0.0234375,-0.0,0.03125,-0.0625,0.03125,0.078125,0.0390625,-0.0546875,-0.0234375,0.0078125,-0.0546875,0.0078125,-0.0546875,0.0546875,0.0078125,-0.046875,0.0390625,-0.109375,-0.03125,-0.0546875,0.0703125,-0.0234375,-0.0234375,0.0625,-0.0078125,-0.015625,0.109375,0.015625,0.015625,-0.0234375,-0.0390625,-0.0390625,-0.1640625,-0.0546875,0.0078125,0.0078125,-0.0625,0.078125,0.0078125,0.03125,-0.015625,-0.0234375,-0.0546875,-0.0390625,0.0625,-0.0625,0.0390625,0.0078125,-0.03125,0.0703125,0.0703125,-0.09375,-0.0078125,-0.046875,0.0546875,-0.015625,-0.078125,0.1953125,-0.0703125,0.078125,-0.0078125,0.078125,-0.1015625,-0.0078125,-0.0859375,0.03125,-0.0703125,-0.0234375,-0.03125,-0.046875,0.0,0.0078125,0.1484375,0.0078125,-0.015625,0.015625,-0.109375,0.0078125,-0.0,0.0078125,-0.078125,-0.046875,0.03125,0.015625,0.0234375,-0.0078125,-0.0,-0.015625,0.046875,-0.0234375,-0.109375,0.0078125,0.2109375,-0.03125,0.0703125,-0.0859375,0.0234375,-0.0390625,0.109375,-0.0,-0.0859375,-0.0078125,-0.0546875,-0.0546875,-0.0390625,0.0625,0.0234375,-0.09375,-0.0,-0.0625,-0.078125,-0.0703125,-0.015625,-0.03125,0.0703125,-0.0,-0.0078125,-0.03125,-0.0390625,0.0703125,0.0703125,0.125,0.109375,-0.0546875,0.015625,-0.0390625,0.125,-0.0234375,0.0078125,-0.09375,0.0,0.0234375,0.125,-0.0,0.0234375,0.078125,-0.09375,0.140625,0.0390625,-0.0,-0.0625,-0.0859375,0.078125,-0.015625,-0.0234375,-0.03125,0.03125,-0.15625,-0.1640625,-0.140625,-0.03125,-0.09375,0.0,0.09375,-0.0078125,-0.09375,-0.015625,0.109375,0.0625,-0.0390625,-0.1796875,0.0859375,0.0625,0.15625,0.1015625,0.015625,-0.03125,0.15625,0.015625,0.09375,0.1328125,0.0546875,0.0390625,-0.046875,0.0625,0.03125,0.1640625,-0.0,0.1015625,0.0234375,0.015625,-0.1015625,-0.109375,0.078125,0.03125,0.1953125,0.078125,0.0234375,0.1796875,0.0078125,0.109375,-0.0078125,0.0546875,-0.0390625,0.046875,-0.0703125,-0.015625,0.1484375,-0.1171875,0.109375,0.0625,-0.0859375,-0.0859375,-0.015625,0.109375,0.0859375,-0.1015625,0.1171875,-0.1015625,-0.140625,-0.078125,-0.078125,0.0703125,0.015625,-0.0078125,0.015625,0.078125,-0.046875,0.1171875,-0.0078125,-0.1328125,-0.078125,-0.0546875,-0.0703125,0.078125,-0.0234375,-0.0390625,-0.1640625,0.1953125,0.078125,-0.0703125,-0.1328125,-0.078125,-0.0859375,-0.0859375,-0.03125,0.0234375,0.0234375,0.0078125,0.0625,-0.046875,-0.03125,-0.046875,-0.078125,-0.0078125,0.0703125,0.09375,0.0546875,-0.0234375,-0.0078125,-0.0,0.0078125,-0.0546875,0.078125,0.0078125,0.0078125,0.015625,0.015625,-0.03125,-0.0,-0.0703125,0.0078125,0.015625,-0.015625,-0.0390625,-0.0,0.0625,-0.03125,0.09375,0.0234375,0.0,0.09375,0.0078125,-0.109375,0.0078125,0.0546875,0.015625,-0.0546875,-0.046875,-0.1640625,-0.0078125,-0.015625,0.0234375,0.0,-0.0234375,0.0625,0.03125,-0.0234375,-0.1015625,-0.015625,0.046875,-0.0703125,-0.0546875,-0.0234375,0.1171875,-0.09375,0.03125,0.0078125,-0.0078125,0.015625,0.0703125,-0.0625,-0.078125,0.015625,0.0,0.0625,0.015625,0.0,0.03125,0.109375,0.015625,-0.0390625,-0.0546875,-0.078125,0.0859375,0.046875,-0.0078125,0.0078125,0.0390625,0.015625,0.03125,0.03125,0.0390625,0.0234375,-0.015625,0.0078125,-0.0390625,0.015625,0.078125,-0.140625,0.015625,-0.125,-0.0078125,-0.03125,0.125,-0.015625,-0.0546875,0.015625,-0.078125,0.0234375,-0.0390625,0.0,0.0078125,0.0703125,-0.015625,0.09375,0.0859375,0.046875,-0.0078125,-0.03125,-0.0390625,-0.0625,0.1015625,0.0703125,-0.0234375,0.015625,-0.046875,0.015625,0.0078125,0.0234375,0.015625,0.1015625,0.0078125,-0.0703125,0.171875,-0.03125,-0.09375,0.03125,0.015625,-0.0234375,-0.015625,-0.0078125,0.0703125,0.0625,-0.03125,0.1171875,-0.0390625,0.03125,-0.1015625,0.0625,0.0390625,0.0,0.03125,0.0234375,-0.015625,0.0703125,0.109375,-0.0234375,-0.0546875,-0.0078125,-0.0546875,0.1640625,0.1171875,-0.078125,0.1875,0.0234375,-0.0390625,-0.046875,0.046875,-0.0078125,0.0,0.03125,-0.203125,0.0625,-0.09375,0.0625,0.0546875,0.03125,-0.0078125,-0.03125,-0.0546875,0.0625,0.1640625,-0.1171875,0.0546875,-0.03125,-0.0390625,0.0078125,0.046875,-0.03125,0.2109375,0.1171875,-0.1171875,-0.0234375,0.03125,0.0546875,0.109375,0.046875,-0.1171875,0.1796875,-0.015625,0.0703125,-0.03125,-0.15625,0.1953125,0.046875,0.0859375,0.109375,0.015625,0.171875,-0.0859375,-0.0390625,0.0,0.0390625,-0.0703125,0.0,-0.015625,0.0859375,0.1484375,0.0703125,0.1328125,-0.140625,0.078125,0.0234375,0.0625,-0.0546875,-0.015625,0.1640625,-0.0625,0.0390625,-0.140625,-0.0546875,0.0546875,0.0078125,0.0390625,-0.0,0.1171875,-0.0546875,-0.078125,-0.0078125,-0.1015625,-0.0703125,-0.0546875,-0.140625,-0.015625,0.0703125,-0.046875,-0.09375,0.03125,-0.1328125,-0.21875,0.015625,0.0234375,0.109375,0.0703125,0.2578125,0.0234375,0.109375,-0.09375,0.1484375,0.0234375,-0.1171875,0.0078125,-0.0078125,0.0,-0.03125,-0.09375,0.0390625,-0.0078125,-0.0703125,-0.0,-0.03125,0.0234375,0.0390625,0.0546875,-0.0703125,0.0625,0.046875,-0.0234375,0.0546875,0.0078125,-0.03125,0.015625,-0.0546875,-0.0625,-0.0859375,-0.0625,-0.0625,-0.0546875,-0.1015625,-0.015625,-0.0078125,0.1875,-0.03125,-0.0546875,0.015625,-0.125,-0.0546875,0.03125,-0.0546875,0.0234375,0.0703125,0.0078125,-0.03125,-0.0,-0.0078125,-0.0234375,-0.0625,-0.046875,0.0078125,0.0390625,0.0,0.046875,0.03125,-0.0390625,-0.03125,-0.1640625,0.046875,0.03125,-0.015625,0.0703125,-0.015625,0.078125,0.09375,-0.1796875,-0.0859375,-0.0390625,-0.0,-0.0546875,-0.0078125,-0.0078125,0.0859375,-0.0390625,0.0546875,-0.0390625,-0.0078125,-0.03125,-0.015625,-0.0234375,0.125,0.0,-0.0234375,0.0078125,-0.015625,-0.0234375,-0.0859375,0.25,0.109375,0.0,-0.0078125,0.0546875,-0.0390625,0.0625,-0.0,-0.0625,0.0078125,0.0234375,-0.0078125,0.0546875,-0.0078125,-0.09375,-0.0078125,0.0,0.0078125,-0.015625,-0.0859375,-0.0390625,-0.0078125,0.0078125,0.03125,0.0078125,-0.046875,-0.0625,-0.0859375,0.0625,-0.0625,0.0234375,0.0546875,-0.0234375,-0.015625,0.046875,0.046875,0.09375,-0.0078125,-0.0390625,0.0,-0.0078125,0.046875,0.0703125,0.0,-0.09375,-0.0078125,0.078125,0.078125,0.0,-0.015625,-0.0234375,0.0078125,0.015625,-0.0703125,-0.03125,-0.0546875,0.015625,0.03125,0.03125,-0.0546875,-0.0390625,0.09375,0.078125,0.0078125,0.0078125,0.0390625,0.0390625,0.0234375,-0.0703125,-0.171875,-0.0078125,-0.0078125,-0.03125,-0.0,0.1328125,-0.03125,0.0859375,-0.109375,-0.0078125,0.1953125,0.0078125,-0.0390625,0.0703125,-0.0234375,-0.0078125,0.0859375,0.0703125,-0.0234375,-0.15625,-0.046875,-0.09375,0.0859375,0.1015625,0.0234375,-0.078125,-0.0234375,0.0546875,0.03125,-0.0703125,0.03125,0.0390625,0.046875,-0.078125,0.0234375,-0.0390625,-0.03125,-0.171875,-0.015625,-0.0234375,-0.1015625,-0.09375,0.03125,0.015625,0.0703125,-0.046875,-0.046875,-0.015625,-0.03125,-0.015625,0.0078125,0.109375,-0.046875,-0.0234375,0.03125,-0.078125,0.015625,-0.0390625,-0.03125,0.2109375,0.0234375,-0.015625,0.0234375,-0.1796875,0.0703125,-0.078125,0.03125,-0.1015625,-0.0859375,0.015625,0.0390625,0.125,-0.09375,-0.0078125,0.0234375,-0.03125,-0.1015625,-0.0234375,-0.0,0.1328125,0.0546875,0.046875,-0.09375,0.0078125,-0.015625,0.0625,0.0390625,0.046875,-0.0546875,-0.09375,0.0234375,-0.0625,0.0,-0.0546875,-0.09375,0.1796875,-0.0703125,-0.078125,-0.0546875,-0.0703125,-0.046875,0.03125,-0.0234375,-0.1015625,-0.015625,-0.015625,0.125,0.1640625,-0.046875,-0.09375,0.078125,0.1484375,-0.03125,0.0703125,-0.0625,-0.0234375,0.0,0.015625,0.0,-0.0,0.078125,-0.0078125,0.0703125,-0.0234375,-0.0,0.0390625,-0.0,0.1171875,-0.03125,0.0703125,-0.0234375,0.0390625,0.0078125,-0.0546875,0.0546875,0.0390625,-0.0625,-0.03125,0.0,-0.0390625,-0.015625,0.078125,0.0703125,0.1171875,0.0,0.015625,-0.0078125,0.015625,0.0078125,-0.0078125,0.046875,-0.015625,0.046875,0.0234375,0.0234375,0.109375,0.015625,-0.0703125,0.03125,0.0390625,0.0625,0.0703125,0.03125,0.109375,0.0,-0.09375,0.0234375,-0.0546875,0.0,-0.09375,0.0390625,-0.0546875,-0.03125,-0.0390625,0.0234375,0.046875,0.0546875,0.0078125,-0.0234375,-0.0859375,0.0859375,-0.046875,-0.1328125,0.015625,0.015625,-0.0859375,-0.0078125,0.0078125,0.0390625,-0.03125,0.0078125,0.0078125,-0.03125,-0.046875,0.0234375,0.0078125,-0.0390625,0.046875,-0.03125,-0.0703125,0.0234375,0.0,-0.0078125,-0.046875,-0.0,0.015625,-0.0,0.109375,0.0,0.0078125,0.0546875,-0.046875,0.0078125,-0.0859375,-0.0625,0.0859375,0.046875,0.0859375,-0.015625,0.0390625,-0.0234375,0.03125,-0.0546875,-0.03125,0.015625,-0.0703125,-0.078125,0.0234375,-0.0546875,-0.03125,-0.046875,-0.0078125,0.078125,-0.046875,0.015625,0.0,0.0234375,-0.015625,-0.0078125,-0.0234375,0.03125,0.015625,0.0,-0.0078125,0.0234375,-0.1484375,-0.15625,0.0078125,-0.0234375,-0.0078125,0.1796875,0.0546875,-0.046875,0.015625,-0.1484375,0.125,0.0078125,0.078125,0.015625,0.0,0.0234375,-0.0546875,0.03125,0.0703125,-0.046875,0.1171875,-0.0234375,0.015625,0.0703125,0.1953125,0.015625,0.03125,-0.0390625,-0.03125,0.09375,-0.0703125,-0.046875,0.1796875,-0.0,-0.125,0.15625,0.0,0.0546875,0.0390625,-0.1640625,0.203125,-0.0,0.0625,0.046875,-0.1171875,-0.1484375,-0.0390625,-0.125,0.1484375,-0.09375,-0.1484375,-0.046875,-0.0234375,-0.125,-0.0546875,0.0234375,-0.15625,-0.109375,0.2890625,0.046875,0.0703125,-0.0625,0.0390625,-0.21875,0.0078125,-0.09375,0.109375,0.171875,0.2109375,0.0703125,-0.140625,-0.0234375,-0.1015625,0.109375,-0.0859375,-0.0234375,0.046875,0.03125,-0.03125,-0.0078125,0.2265625,0.0859375,-0.015625,0.015625,0.0,-0.1171875,0.1640625,0.171875,0.1953125,-0.03125,-0.0078125,0.0859375,-0.0078125,0.03125,-0.0078125,0.109375,0.0546875,-0.0,0.125,-0.1015625,-0.03125,0.171875,-0.0,-0.1796875,0.1484375,-0.1015625,-0.125,0.109375,0.015625,0.0625,0.1328125,-0.03125,0.0703125,0.140625,0.03125,0.0625,-0.0703125,-0.125,-0.015625,-0.0,-0.078125,0.1875,0.1171875,0.0078125,-0.1875,0.1796875,-0.109375,-0.1328125,0.03125,0.03125,-0.015625,-0.03125,-0.015625,0.0,0.0078125,-0.015625,0.109375,-0.0078125,0.0,-0.0234375,0.0078125,-0.0625,-0.0,0.0,-0.0234375,-0.03125,-0.0078125,-0.046875,-0.03125,-0.0234375,-0.0390625,-0.0078125,-0.0703125,-0.015625,-0.03125,-0.015625,-0.0234375,-0.0625,-0.0078125,0.015625,-0.0546875,0.015625,0.0859375,-0.078125,0.046875,0.03125,-0.1171875,0.0078125,-0.0234375,-0.046875,0.015625,-0.0546875,0.0390625,-0.03125,-0.0859375,-0.03125,-0.125,0.1328125,-0.0390625,-0.0390625,0.0390625,-0.015625,0.0078125,0.0234375,-0.015625,-0.0703125,0.0703125,0.0078125,-0.015625,0.0234375,0.046875,-0.0703125,0.0390625,0.0546875,0.0,-0.0859375,-0.0078125,-0.015625,-0.0234375,0.1015625,-0.046875,0.0,-0.0390625,-0.0546875,-0.03125,-0.0078125,-0.0,0.078125,0.015625,-0.0,-0.03125,-0.078125,0.03125,0.0,0.015625,-0.046875,-0.03125,-0.0390625,-0.046875,0.0,-0.0,0.046875,0.0859375,-0.046875,-0.046875,-0.0859375,-0.0859375,-0.0625,-0.015625,-0.0546875,-0.1171875,0.09375,0.1484375,0.0078125,0.0703125,0.0078125,-0.015625,0.015625,-0.015625,0.0390625,0.0390625,-0.0,-0.0078125,-0.0390625,0.015625,-0.0078125,-0.0,-0.015625,-0.046875,-0.0078125,0.0234375,-0.0703125,-0.0234375,0.078125,-0.0078125,-0.0703125,-0.015625,-0.0390625,0.0546875,-0.0625,0.03125,-0.078125,-0.0546875,0.140625,0.046875,0.0078125,0.03125,0.0859375,-0.03125,0.0625,-0.046875,-0.0703125,0.0078125,0.015625,-0.078125,-0.0625,0.015625,-0.0625,-0.0390625,0.0234375,0.0,0.0703125,-0.046875,0.09375,-0.03125,-0.0703125,-0.1796875,-0.015625,-0.0546875,0.03125,0.0,0.171875,-0.0546875,-0.0390625,0.1328125,0.015625,0.0078125,0.0859375,0.0625,0.1015625,-0.0625,-0.03125,0.046875,-0.0390625,0.0078125,0.0234375,0.0703125,0.0078125,0.125,-0.015625,0.09375,0.0234375,-0.0625,0.1015625,-0.0859375,-0.109375,0.0390625,0.171875,-0.0625,0.0234375,0.03125,0.0546875,-0.0625,-0.1953125,-0.0703125,0.1015625,0.015625,-0.0,-0.0078125,-0.015625,-0.09375,0.0078125,0.0625,-0.015625,-0.03125,-0.0,0.015625,0.03125,0.015625,0.03125,0.078125,0.0625,0.078125,0.0,0.1796875,-0.0390625,-0.0625,0.1015625,-0.0703125,-0.046875,0.1171875,0.015625,-0.0546875,-0.015625,0.15625,-0.109375,-0.0234375,-0.046875,0.0546875,-0.0546875,-0.078125,-0.109375,0.0859375,0.0234375,-0.015625,-0.0390625,-0.1015625,0.0,-0.046875,0.0546875,0.1640625,0.1171875,0.03125,-0.0234375,-0.015625,0.0390625,-0.0,-0.109375,0.0546875,-0.0390625,0.0,0.0703125,-0.09375,0.015625,0.0234375,0.0234375,0.0078125,0.0,0.015625,-0.046875,-0.0,0.0,0.0390625,-0.0390625,0.15625,-0.0234375,0.046875,0.0078125,-0.0234375,0.0078125,0.09375,-0.0625,-0.0859375,0.046875,0.109375,-0.1328125,0.0703125,-0.0390625,-0.0234375,0.0234375,-0.0234375,-0.015625,-0.0390625,-0.03125,-0.0078125,0.015625,0.0546875,-0.0078125,0.015625,-0.0859375,0.078125,-0.0234375,-0.0078125,-0.0625,0.0546875,-0.0703125,-0.0390625,-0.1015625,-0.0703125,0.0078125,0.0390625,0.0078125,-0.0859375,-0.0546875,0.0078125,-0.109375,-0.109375,0.0,0.0078125,-0.0234375,-0.0546875,0.09375,0.0234375,-0.0859375,0.0078125,0.0078125,-0.015625,0.0546875,-0.03125,-0.015625,0.0078125,0.0546875,-0.1171875,0.03125,-0.0234375,0.0625,-0.0078125,-0.0,0.0625,0.0078125,-0.0,0.0078125,0.015625,0.0234375,-0.0,-0.109375,0.125,0.0234375,0.03125,-0.015625,0.0234375,-0.015625,-0.0390625,0.0546875,-0.015625,-0.015625,0.0,-0.0625,-0.0078125,0.0,-0.09375,-0.0703125,0.0703125,-0.1640625,-0.0078125,-0.0234375,0.046875,-0.0390625,0.1953125,0.0078125,0.1640625,0.015625,-0.1484375,-0.0078125,0.0546875,-0.015625,-0.0234375,0.078125,-0.1484375,-0.0390625,0.0234375,0.0703125,-0.015625,0.015625,-0.0234375,0.0,0.046875,0.0234375,-0.0625,0.0625,-0.0234375,0.03125,-0.03125,-0.0390625,0.0625,0.03125,-0.0,0.0234375,0.1640625,0.171875,0.046875,-0.0390625,-0.0625,0.0703125,-0.03125,-0.0546875,0.0078125,-0.015625,0.046875,0.1640625,0.0234375,0.21875,0.0390625,-0.09375,0.03125,0.1015625,0.0078125,0.046875,-0.0390625,-0.1328125,-0.046875,0.0546875,-0.1328125,-0.09375,0.0234375,0.0859375,-0.0078125,0.015625,-0.0234375,-0.15625,-0.0390625,-0.015625,-0.09375,0.140625,-0.0234375,-0.078125,0.0078125,-0.140625,-0.09375,0.015625,0.0546875,0.078125,0.1328125,0.0,-0.0234375,-0.015625,0.0625,0.0546875,-0.0390625,0.203125,-0.0546875,-0.1015625,-0.0390625,0.0078125,-0.015625,-0.015625,-0.046875,0.1015625,0.0078125,-0.0078125,-0.0625,0.015625,-0.0078125,-0.015625,-0.015625,-0.09375,-0.0390625,0.046875,-0.0546875,-0.078125,-0.0234375,0.1015625,-0.0625,0.0,-0.046875,-0.0078125,0.046875,-0.140625,-0.0390625,-0.1015625,0.03125,-0.0078125,0.0234375,0.3046875,-0.0703125,-0.0078125,0.0546875,0.0078125,0.0625,0.0,0.1484375,-0.03125,-0.1484375,-0.0078125,0.015625,0.0859375,-0.0625,0.0390625,-0.046875,0.0078125,-0.078125,-0.046875,-0.1015625,0.078125,0.0625,-0.125,0.09375,-0.0546875,0.0390625,0.0078125,-0.03125,0.0546875,-0.015625,0.0625,0.078125,0.0234375,0.140625,-0.0,-0.09375,-0.078125,0.015625,0.1171875,0.0,-0.0234375,0.0078125,-0.046875,-0.015625,0.0078125,-0.0625,-0.0078125,0.0078125,-0.046875,0.0625,0.0703125,-0.0078125,-0.0,-0.0625,0.0,-0.0078125,-0.109375,-0.09375,-0.0390625,0.03125,0.03125,0.03125,-0.03125,0.0234375,-0.03125,0.0390625,0.0625,-0.015625,-0.0,0.125,-0.015625,-0.0390625,0.015625,-0.0703125,-0.0078125,0.1328125,-0.0,-0.0390625,0.21875,-0.015625,0.21875,0.1328125,0.1171875,0.03125,0.0078125,0.0234375,-0.0,0.0078125,0.015625,0.0625,0.0,-0.03125,0.15625,-0.0390625,-0.03125,-0.015625,-0.03125,0.09375,0.0078125,-0.078125,0.0703125,0.0078125,-0.0078125,0.03125,-0.03125,-0.0625,0.0546875,0.0546875,0.03125,-0.09375,-0.015625,0.015625,0.03125,0.078125,-0.0,0.1328125,-0.078125,-0.0078125,0.0859375,0.0,-0.078125,0.0625,-0.0,0.0546875,0.09375,-0.0234375,0.015625,0.015625,-0.0,-0.0078125,-0.015625,-0.0234375,-0.0625,0.0546875,0.1171875,0.0625,-0.0,0.015625,0.0703125,-0.0234375,0.0078125,-0.0,-0.0078125,-0.09375,0.0078125,-0.0,-0.015625,-0.03125,0.0390625,0.0078125,-0.078125,0.03125,0.0703125,-0.0859375,-0.0390625,0.015625,-0.0234375,0.0390625,0.015625,0.015625,-0.046875,0.046875,-0.015625,0.0390625,-0.0078125,-0.0,0.0234375,-0.109375,-0.015625,-0.0390625,-0.0859375,0.03125,0.0234375,0.125,-0.03125,-0.109375,-0.0546875,0.0703125,0.0234375,0.03125,-0.015625,-0.0859375,-0.015625,0.0390625,0.1015625,-0.0625,-0.03125,0.0703125,-0.0625,0.0390625,0.03125,0.046875,-0.1640625,0.046875,-0.0078125,0.03125,0.0,-0.0625,-0.0546875,0.0625,0.0078125,-0.03125,-0.0234375,-0.046875,0.109375,0.109375,0.0859375,-0.0703125,-0.03125,0.0625,0.0703125,-0.0,0.109375,0.09375,-0.015625,-0.03125,0.1640625,0.0859375,-0.0703125,-0.0703125,-0.0234375,-0.03125,0.0234375,0.0,0.1171875,-0.03125,-0.1015625,-0.0625,-0.078125,0.078125,-0.0234375,0.0,0.0234375,0.0234375,0.0546875,-0.0234375,-0.03125,0.0234375,-0.0234375,0.0546875,0.0625,0.0078125,0.0546875,-0.0703125,0.0078125,-0.0234375,-0.0234375,-0.0390625,-0.046875,0.046875,-0.015625,0.0859375,-0.0546875,-0.03125,-0.015625,-0.1015625,-0.0859375,0.0625,-0.015625,-0.15625,-0.1484375,0.015625,0.109375,-0.1171875,-0.015625,0.1796875,-0.0234375,-0.0546875,-0.046875,-0.0078125,-0.0546875,-0.09375,0.0234375,-0.078125,-0.0234375,-0.078125,0.171875,-0.0,-0.0703125,0.015625,-0.0078125,0.0078125,-0.046875,-0.0625,-0.0,0.015625,-0.0703125,-0.0234375,0.09375,0.046875,-0.015625,0.0078125,0.0625,-0.015625,-0.0078125,0.0625,-0.0625,0.0,-0.0,-0.0703125,-0.0078125,0.0234375,0.046875,0.0703125,0.015625,0.0234375,0.109375,0.0234375,0.0078125,-0.015625,0.0703125,-0.0859375,-0.0390625,0.1328125,-0.140625,-0.0234375,0.03125,0.03125,-0.0390625,-0.0078125,0.03125,0.0078125,-0.0,0.0390625,0.0078125,-0.0390625,-0.015625,-0.0546875,0.046875,0.078125,-0.0703125,0.0078125,0.078125,0.0859375,0.0546875,-0.0625,0.0,-0.03125,0.03125,-0.03125,-0.0234375,0.0703125,0.0390625,0.03125,-0.0234375,-0.0078125,0.015625,-0.0546875,-0.0234375,0.0,-0.015625,-0.015625,-0.0234375,0.0078125,0.0234375,0.0,0.0546875,-0.0,0.0078125,0.015625,0.0546875,0.0,0.0390625,-0.015625,0.09375,-0.015625,0.0078125,0.015625,-0.0,0.0859375,-0.0390625,-0.015625,-0.03125,-0.015625,-0.09375,0.0078125,0.1796875,-0.0390625,-0.0,0.09375,0.0390625,0.140625,-0.0390625,0.0234375,-0.0,-0.0,-0.078125,0.0,0.0078125,-0.09375,0.015625,-0.078125,0.0625,-0.0546875,-0.0703125,-0.0703125,-0.03125,-0.015625,0.0234375,-0.03125,0.0,0.0390625,0.015625,-0.0546875,-0.0703125,0.015625,0.0859375,-0.0390625,0.03125,0.0625,-0.0,-0.0078125,0.0546875,0.03125,0.0078125,-0.0,-0.078125,-0.0078125,-0.015625,0.0859375,-0.1640625,0.03125,0.0234375,0.109375,-0.0546875,0.1484375,0.0078125,0.1328125,0.140625,-0.1015625,-0.0078125,0.0703125,-0.1171875,-0.125,0.09375,-0.0703125,-0.09375,0.1015625,0.0234375,-0.0546875,-0.03125,0.0546875,0.1640625,0.0625,0.1484375,-0.125,-0.0703125,-0.078125,-0.09375,-0.046875,0.078125,-0.015625,-0.046875,0.046875,-0.0,-0.015625,-0.046875,-0.0390625,0.078125,-0.140625,0.0859375,-0.0390625,-0.046875,0.234375,-0.1484375,0.0390625,-0.046875,0.03125,-0.171875,0.0625,-0.109375,0.1640625,0.0546875,-0.0546875,-0.0703125,-0.2109375,0.0,0.1953125,-0.0625,0.1640625,0.03125,0.015625,0.125,0.1640625,-0.0,0.0078125,0.0625,-0.0546875,0.0234375,0.015625,0.046875,0.109375,0.0234375,-0.09375,-0.0078125,-0.0859375,0.0390625,0.1015625,-0.0703125,-0.015625,0.1015625,0.0703125,0.0859375,-0.0078125,0.0078125,-0.140625,-0.1015625,-0.0546875,-0.0390625,0.03125,0.21875,-0.0703125,-0.0546875,-0.0390625,-0.046875,-0.03125,0.1484375,-0.0703125,0.0625,-0.078125,-0.0,-0.0625,0.09375,-0.0703125,0.0234375,0.109375,-0.015625,0.0625,-0.0234375,0.0390625,-0.109375,0.0390625,0.09375,-0.125,-0.0390625,-0.0390625,-0.015625,-0.09375,-0.03125,0.15625,0.1328125,-0.0078125,0.0859375,-0.109375,0.015625,-0.0546875,-0.140625,-0.09375,0.0390625,-0.046875,-0.0078125,0.0078125,-0.0078125,-0.0,0.0078125,0.046875,0.0390625,0.0390625,0.0390625,-0.03125,0.0859375,-0.0078125,0.015625,0.0390625,-0.0078125,-0.0546875,0.0625,0.1015625,-0.0234375,0.0625,0.0234375,0.03125,-0.0546875,0.0390625,-0.03125,0.0234375,-0.015625,0.0234375,0.0625,-0.0234375,-0.0546875,0.015625,-0.015625,0.0234375,-0.0,-0.1328125,0.0390625,0.1328125,0.03125,0.0,-0.0234375,-0.046875,-0.0390625,0.0390625,0.015625,0.0625,0.0078125,0.1328125,0.0546875,-0.0546875,0.015625,0.0,-0.0078125,-0.0234375,-0.078125,0.03125,-0.03125,-0.0625,0.0859375,-0.0546875,-0.015625,0.0625,-0.0546875,0.0703125,-0.0078125,0.015625,0.0625,0.046875,-0.0,-0.015625,-0.03125,0.09375,-0.0,0.015625,0.0703125,0.0078125,0.0,-0.0703125,0.015625,0.0234375,-0.0546875,-0.09375,0.03125,0.0625,-0.0,-0.1171875,-0.078125,-0.0078125,0.0234375,0.1015625,0.0234375,-0.0,0.078125,-0.0390625,0.078125,-0.09375,0.046875,-0.03125,0.1484375,0.0,-0.0703125,-0.015625,0.0390625,-0.140625,-0.046875,0.0234375,0.0078125,0.0234375,-0.015625,0.0546875,0.0,0.0078125,-0.0234375,0.125,0.015625,0.0078125,0.0,0.0234375,0.046875,0.0546875,0.0078125,-0.0234375,0.046875,0.0078125,-0.0,0.015625,0.1875,0.0078125,-0.046875,0.046875,0.0,0.0234375,0.0234375,0.1484375,0.125,-0.0390625,0.0,0.046875,0.015625,0.171875,0.0546875,0.015625,0.140625,-0.046875,0.1875,0.0234375,0.078125,-0.0390625,0.0859375,-0.0390625,-0.09375,-0.0703125,-0.1875,-0.0390625,-0.1953125,0.0625,-0.046875,-0.0703125,-0.0546875,-0.0,0.0078125,-0.0546875,-0.0859375,-0.078125,0.0234375,0.015625,0.0078125,-0.046875,-0.015625,0.0,-0.03125,-0.15625,-0.0859375,-0.0078125,-0.0390625,-0.0234375,-0.0,-0.0078125,0.09375,-0.078125,-0.0,-0.1171875,-0.0859375,0.0703125,-0.140625,-0.1953125,0.0546875,-0.1015625,0.0703125,-0.09375,0.0859375,0.3125,0.109375,0.1171875,-0.0078125,0.078125,0.0546875,0.0078125,-0.0078125,-0.125,-0.0078125,0.1015625,-0.0703125,-0.0390625,0.0546875,-0.0234375,0.0078125,-0.15625,-0.046875,0.265625,0.0234375,-0.078125,-0.1015625,-0.078125,-0.03125,-0.0859375,0.015625,-0.0625,-0.015625,-0.078125,-0.0625,0.1171875,0.0703125,0.1640625,0.046875,0.15625,0.15625,0.0703125,-0.09375,-0.0234375,-0.0,0.03125,0.03125,0.0625,0.09375,0.015625,0.0234375,0.15625,0.015625,0.0078125,0.0234375,0.203125,0.078125,0.109375,-0.1796875,0.046875,0.0703125,-0.1640625,-0.0234375,0.0703125,0.0390625,0.171875,0.109375,-0.0625,-0.0390625,0.015625,0.0234375,-0.046875,-0.0,0.0078125,-0.0,0.03125,-0.0,-0.046875,-0.015625,0.0234375,-0.0,-0.0390625,0.1015625,-0.0234375,0.0078125,0.046875,-0.03125,-0.0234375,0.0546875,0.0859375,-0.015625,0.0,-0.0234375,0.1171875,0.0859375,-0.015625,0.0078125,-0.015625,-0.078125,-0.0390625,-0.015625,0.046875,0.0,-0.0390625,0.0078125,-0.0078125,-0.0,0.0390625,-0.0,0.015625,0.0234375,-0.03125,0.09375,-0.0703125,0.015625,0.0546875,0.0078125,0.109375,0.015625,0.0625,0.046875,-0.0859375,-0.015625,0.0078125,0.078125,-0.0546875,0.1171875,-0.09375,0.046875,0.109375,-0.015625,-0.0234375,-0.046875,0.015625,-0.0390625,-0.0234375,0.0859375,-0.0546875,0.03125,-0.03125,0.015625,0.125,0.0390625,0.015625,0.1171875,0.0,-0.0234375,0.1015625,0.015625,0.0078125,-0.0859375,0.046875,0.0703125,-0.03125,-0.0,0.0,0.0546875,-0.0234375,0.0234375,0.03125,0.0234375,0.0,0.0703125,-0.03125,0.0078125,-0.1015625,0.0859375,-0.09375,0.0390625,-0.0390625,0.0390625,0.109375,0.0234375,0.0390625,-0.0078125,0.0703125,0.0234375,-0.09375,0.0078125,0.0859375,0.0703125,-0.1171875,0.0703125,-0.0390625,0.0546875,0.0625,0.0234375,0.0078125,0.0546875,0.03125,-0.0,0.0625,0.03125,-0.046875,-0.0390625,0.0078125,0.1953125,0.0390625,-0.03125,-0.1328125,-0.109375,-0.0,0.0078125,-0.03125,0.046875,0.0703125,0.0,-0.0859375,0.0859375,0.2109375,0.015625,0.0546875,-0.0703125,-0.1484375,-0.0703125,-0.0078125,-0.0625,-0.0234375,-0.015625,0.1328125,0.0078125,0.0546875,-0.0078125,0.2734375,-0.0078125,-0.015625,-0.0703125,-0.0078125,-0.0546875,0.0390625,-0.0,0.0,0.0625,0.1796875,-0.1015625,0.078125,-0.09375,0.0625,0.1640625,-0.0625,-0.0625,-0.0625,-0.109375,-0.0625,0.0234375,0.0078125,0.0078125,0.046875,0.0078125,-0.15625,0.0546875,-0.0546875,-0.0625,-0.078125,-0.0859375,0.0,-0.125,0.046875,-0.1640625,-0.0234375,-0.125,-0.03125,0.1171875,0.09375,-0.0078125,0.0625,0.0234375,-0.109375,-0.0234375,-0.015625,-0.0546875,-0.0546875,-0.1640625,-0.1015625,0.0546875,0.078125,0.09375,0.078125,0.078125,0.0234375,-0.1796875,0.1015625,0.0078125,0.0546875,-0.0546875,-0.078125,0.1171875,0.0234375,0.0078125,-0.03125,0.0234375,-0.0625,-0.0,-0.0234375,-0.03125,0.078125,0.0625,-0.015625,0.0703125,0.0390625,0.109375,0.03125,0.078125,-0.0390625,-0.03125,0.1015625,-0.109375,0.09375,0.125,0.046875,-0.2109375,0.109375,-0.2109375,0.015625,0.1171875,-0.0703125,0.0546875,-0.1484375,-0.0078125,-0.09375,-0.0390625,0.046875,-0.03125,-0.0078125,0.0078125,0.0546875,-0.0390625,-0.015625,-0.0,0.0078125,-0.0078125,-0.0,-0.0,-0.03125,-0.03125,-0.0625,-0.0078125,0.0078125,-0.0703125,0.015625,-0.0078125,0.0859375,-0.0234375,0.0390625,0.0078125,0.0546875,0.046875,0.0234375,-0.046875,0.0390625,0.046875,-0.03125,0.0078125,0.0234375,0.0,-0.0390625,0.0,0.046875,0.0390625,-0.0078125,-0.0234375,-0.078125,0.015625,0.0703125,-0.0,-0.0625,0.0078125,-0.0859375,0.0,0.015625,0.1171875,0.1640625,0.03125,-0.015625,-0.0625,-0.015625,0.046875,-0.0234375,0.0,0.078125,0.1484375,0.015625,0.0234375,-0.1015625,0.046875,-0.046875,-0.03125,0.0,0.1171875,0.0078125,-0.0390625,0.015625,-0.046875,-0.0234375,-0.046875,0.109375,-0.03125,0.1171875,0.0234375,0.0234375,-0.0390625,0.015625,-0.03125,-0.015625,0.0078125,0.03125,0.0,-0.015625,0.015625,0.015625,0.0,-0.0390625,0.0,0.0,0.0078125,-0.0078125,0.0078125,0.0234375,0.0625,-0.0234375,0.15625,-0.015625,-0.0,0.0859375,0.0234375,0.0078125,0.0390625,0.0625,-0.0234375,-0.0078125,-0.015625,0.0,-0.015625,-0.0625,-0.015625,0.0390625,0.046875,-0.0234375,-0.0390625,-0.078125,-0.0546875,-0.046875,0.046875,-0.0,0.046875,0.015625,-0.0078125,-0.0390625,0.1015625,0.0078125,-0.0625,0.015625,0.1484375,-0.1640625,-0.1015625,-0.0859375,0.03125,0.109375,-0.078125,0.21875,-0.0625,-0.1015625,0.2109375,-0.015625,-0.0859375,0.0234375,-0.0078125,-0.0625,0.015625,-0.0,-0.1015625,0.1015625,-0.078125,0.125,-0.0859375,-0.03125,-0.03125,-0.1328125,-0.0625,-0.0546875,-0.046875,-0.0625,0.0625,-0.0625,0.0078125,-0.0625,-0.0546875,-0.0078125,0.1171875,0.09375,0.0703125,-0.0546875,-0.046875,0.0390625,-0.0234375,0.0,0.0234375,-0.0859375,0.015625,-0.046875,-0.0390625,0.1171875,-0.0703125,-0.0390625,-0.0390625,0.015625,0.0546875,0.2109375,0.0859375,-0.0625,-0.1171875,-0.0546875,-0.0625,-0.1953125,-0.078125,0.015625,-0.0625,-0.0859375,0.0,-0.0703125,-0.078125,0.046875,-0.0625,0.1328125,0.015625,-0.1171875,-0.0078125,-0.0703125,0.09375,-0.0390625,0.03125,0.046875,-0.078125,-0.0703125,0.0390625,0.0546875,0.0625,0.015625,-0.0234375,-0.03125,-0.140625,-0.078125,-0.125,-0.0078125,-0.015625,0.1171875,0.09375,-0.0078125,0.015625,0.09375,0.015625,0.015625,-0.0234375,-0.0859375,-0.09375,0.2421875,0.0234375,-0.046875,-0.0859375,0.0078125,0.0078125,0.046875,-0.078125,-0.0,-0.1484375,0.1640625,-0.1328125,0.0859375,-0.0234375,-0.015625,-0.015625,0.125,-0.03125,-0.0703125,-0.1640625,-0.0625,0.109375,-0.078125,-0.0546875,-0.0390625,-0.0,-0.0234375,0.015625,-0.046875,0.0234375,0.0078125,0.0390625,0.03125,-0.0390625,0.078125,0.0078125,0.03125,0.0234375,-0.0234375,0.0234375,0.015625,0.015625,0.0859375,0.03125,-0.0234375,-0.03125,0.0234375,0.0234375,0.03125,0.0703125,0.0390625,-0.0,0.015625,0.0234375,-0.015625,-0.0390625,-0.0234375,-0.015625,-0.0703125,0.0,0.0,0.046875,-0.0078125,-0.0234375,-0.0625,-0.0078125,0.0,-0.015625,0.0625,-0.03125,0.1171875,-0.03125,0.0703125,0.0703125,-0.03125,0.0546875,-0.0625,-0.015625,-0.0,0.0,-0.0078125,-0.0390625,0.03125,-0.0546875,-0.015625,-0.0390625,0.0078125,-0.0234375,0.0703125,0.140625,-0.0,-0.0234375,-0.0078125,-0.015625,-0.0078125,0.0234375,-0.0390625,-0.03125,0.015625,0.0078125,0.0703125,0.1015625,-0.03125,0.0078125,0.0390625,-0.0703125,-0.0078125,-0.078125,-0.0390625,-0.015625,-0.0078125,0.015625,0.0234375,-0.0,-0.03125,0.046875,0.03125,0.0078125,-0.0078125,0.0078125,-0.03125,0.09375,0.0078125,-0.03125,0.1953125,0.0546875,0.078125,-0.0390625,0.015625,0.015625,0.0234375,0.0234375,-0.0078125,0.015625,-0.0546875,0.0234375,0.03125,-0.03125,-0.0234375,-0.0234375,0.03125,0.03125,0.046875,0.015625,0.015625,0.046875,-0.0546875,-0.0078125,0.09375,0.0,-0.0,0.0625,-0.140625,-0.1875,-0.0078125,0.0390625,-0.046875,-0.0078125,-0.0078125,0.0546875,-0.0625,-0.015625,0.09375,0.0390625,-0.203125,0.0625,-0.0078125,-0.0078125,0.0234375,-0.0625,-0.09375,-0.015625,0.0078125,0.0234375,-0.0625,0.0,0.15625,0.046875,0.0625,0.0390625,0.21875,0.1953125,-0.015625,-0.0859375,0.0390625,0.0234375,0.1484375,0.078125,0.015625,-0.046875,0.0234375,0.1171875,0.0703125,-0.1484375,-0.09375,-0.0859375,0.0546875,-0.03125,-0.0859375,-0.03125,-0.03125,0.015625,0.0078125,-0.0078125,-0.0234375,0.0,-0.1953125,-0.125,-0.1484375,-0.015625,0.09375,0.0703125,0.0859375,0.0546875,0.046875,-0.1171875,0.09375,-0.1015625,-0.09375,-0.0625,0.015625,0.1015625,0.1484375,0.078125,0.078125,0.0703125,0.03125,-0.0078125,-0.0390625,-0.0703125,0.1171875,-0.1171875,0.1015625,0.0859375,0.125,0.0859375,-0.109375,-0.0625,0.0703125,0.0234375,0.0859375,-0.015625,0.125,0.0,0.0625,-0.046875,0.0234375,-0.0625,-0.1171875,-0.09375,-0.0703125,0.03125,0.0859375,0.046875,-0.109375,-0.1875,-0.046875,-0.234375,-0.0,0.03125,0.078125,-0.0390625,0.15625,0.203125,0.1328125,0.1171875,-0.1640625,0.0703125,0.015625,-0.140625,0.0625,0.1015625,0.0703125,-0.015625,-0.046875,-0.0703125,0.171875,0.046875,0.015625,-0.0078125,-0.046875];

weight_1x1 = [-0.015625,0.0390625,-0.0078125,0.0,0.0078125,-0.0078125,-0.0078125,-0.0546875,-0.0546875,-0.015625,-0.0078125,-0.0234375,-0.0234375,-0.015625,0.015625,0.109375,0.0,0.0,0.0078125,-0.0078125,0.015625,0.0078125,0.0234375,-0.0078125,0.0,-0.046875,-0.046875,-0.0234375,-0.015625,-0.0234375,0.0234375,-0.03125,-0.0546875,-0.0,0.03125,0.046875,-0.0234375,-0.0078125,-0.0234375,-0.0234375,-0.046875,0.0234375,-0.03125,0.0234375,-0.0546875,-0.0234375,-0.0546875,-0.0234375,0.03125,0.0234375,-0.0078125,-0.0,-0.0234375,0.0703125,0.0234375,-0.015625,0.0078125,-0.046875,-0.0234375,0.0,-0.03125,0.0390625,0.0234375,-0.015625,-0.0546875,0.03125,0.046875,-0.046875,-0.0625,0.0078125,0.0859375,-0.0078125,0.0625,-0.015625,0.171875,0.0,-0.015625,-0.03125,0.046875,0.171875,-0.015625,-0.0625,0.03125,0.0859375,0.046875,-0.0390625,0.0234375,-0.0234375,-0.03125,0.0234375,-0.0546875,-0.0703125,-0.046875,-0.015625,-0.015625,0.015625,0.0078125,0.0234375,0.1015625,0.0703125,-0.0234375,0.0234375,0.109375,-0.0625,-0.0859375,-0.0703125,-0.046875,-0.046875,-0.046875,0.03125,-0.0546875,0.03125,-0.0,-0.015625,0.03125,0.03125,-0.0390625,-0.03125,0.125,0.0234375,-0.0390625,-0.046875,0.015625,-0.03125,-0.046875,0.0,0.015625,0.046875,-0.0078125,-0.03125,0.0,-0.046875,0.109375,-0.03125,0.0703125,-0.078125,0.0703125,0.0078125,-0.078125,0.03125,0.0390625,0.0078125,-0.078125,0.0078125,-0.015625,0.0,-0.03125,-0.0546875,0.0234375,-0.0625,0.0078125,-0.0546875,-0.0234375,-0.0859375,-0.03125,0.0234375,0.015625,-0.0625,0.0625,-0.078125,-0.0078125,0.015625,-0.09375,-0.046875,0.0625,0.03125,-0.03125,0.0859375,-0.0078125,-0.0703125,0.0234375,0.046875,0.03125,-0.0078125,0.0234375,0.046875,0.0,-0.0,0.015625,0.03125,0.03125,-0.03125,-0.015625,-0.0703125,0.0625,0.125,0.03125,0.0625,0.0546875,-0.03125,0.0234375,-0.0078125,-0.0078125,-0.015625,0.0390625,-0.03125,-0.03125,-0.0078125,-0.0,0.015625,0.0078125,-0.0234375,-0.0234375,-0.0078125,-0.0234375,0.03125,-0.03125,-0.015625,0.03125,-0.0234375,-0.03125,-0.03125,-0.0234375,0.015625,-0.0078125,-0.03125,0.0078125,0.0390625,0.0078125,-0.0078125,-0.015625,-0.03125,0.0234375,0.0,-0.015625,0.0078125,-0.0703125,0.046875,-0.015625,0.03125,-0.0078125,-0.0234375,-0.0859375,-0.03125,0.0078125,-0.0703125,-0.0390625,-0.0234375,0.0078125,-0.0625,-0.0078125,0.03125,0.0390625,-0.0234375,0.0234375,0.0234375,0.03125,-0.0234375,-0.0703125,-0.078125,0.1328125,-0.1171875,0.0234375,0.1484375,0.0234375,-0.0078125,-0.0390625,0.046875,-0.078125,0.0625,0.1015625,-0.0234375,-0.0078125,0.03125,0.0546875,-0.046875,0.0390625,-0.0078125,0.015625,-0.03125,0.0,-0.0078125,0.015625,-0.0234375,0.0234375,-0.015625,-0.03125,-0.0859375,-0.0546875,-0.0078125,0.0390625,0.0703125,-0.1015625,-0.0234375,0.03125,-0.015625,0.046875,-0.0625,-0.046875,-0.0,-0.0234375,-0.0625,-0.0625,0.0,0.0859375,-0.0390625,-0.015625,-0.015625,0.0390625,-0.0390625,0.0078125,0.0390625,-0.0546875,-0.0234375,0.03125,-0.0078125,-0.0,-0.0390625,0.015625,-0.0078125,0.0390625,-0.0390625,-0.0078125,0.015625,-0.015625,-0.0625,-0.0078125,-0.0,0.0703125,0.046875,-0.015625,0.015625,-0.015625,0.03125,-0.046875,-0.015625,0.0625,0.0078125,0.0703125,-0.0,-0.0078125,0.0078125,-0.015625,-0.0078125,0.03125,-0.0546875,0.0078125,0.03125,0.0,0.0546875,-0.03125,-0.015625,0.0234375,-0.046875,0.015625,-0.0078125,-0.046875,-0.03125,-0.0078125,-0.015625,-0.0234375,0.0078125,0.046875,0.0234375,-0.015625,-0.015625,0.0546875,-0.0078125,-0.015625,0.015625,0.0390625,-0.03125,0.0078125,-0.015625,0.03125,-0.03125,-0.0390625,-0.0078125,0.0234375,0.0625,-0.0390625,0.015625,-0.03125,0.0234375,0.0078125,-0.078125,0.0703125,-0.0,0.0,-0.0078125,-0.0078125,-0.0234375,-0.0234375,0.015625,0.0390625,0.0078125,-0.0078125,-0.0546875,-0.0234375,0.0234375,-0.0390625,-0.0,0.03125,0.015625,0.046875,0.0234375,0.015625,0.0546875,0.015625,-0.015625,0.0234375,-0.015625,-0.03125,-0.0234375,0.0078125,0.0078125,0.0234375,0.0390625,-0.03125,0.015625,-0.046875,0.0390625,-0.0078125,-0.0625,-0.0234375,-0.0390625,-0.0078125,-0.0078125,-0.0546875,0.015625,-0.0,-0.03125,0.015625,-0.03125,0.0625,0.015625,0.046875,-0.015625,0.0390625,0.0078125,-0.0,-0.078125,0.0078125,-0.015625,-0.078125,0.015625,-0.046875,0.0078125,-0.0234375,-0.0546875,-0.0234375,-0.0078125,-0.0234375,0.03125,0.046875,-0.015625,-0.0234375,-0.0078125,0.015625,0.0078125,0.015625,0.046875,-0.046875,0.0,-0.0390625,0.0625,-0.0625,0.0078125,-0.015625,0.0625,-0.0625,0.03125,0.0234375,-0.0625,-0.0390625,-0.078125,-0.0546875,-0.0390625,-0.0625,-0.0078125,-0.0390625,-0.0,-0.046875,0.15625,-0.0,0.0703125,0.03125,0.1171875,-0.0625,0.140625,-0.0,-0.0234375,0.0390625,0.046875,-0.109375,0.03125,-0.0078125,-0.03125,0.1484375,0.046875,-0.046875,-0.0234375,0.0390625,-0.0390625,0.0546875,0.03125,-0.0234375,-0.0234375,-0.0,-0.03125,-0.015625,-0.09375,-0.0234375,-0.1015625,-0.046875,-0.0234375,-0.0390625,0.078125,-0.0078125,0.0078125,0.0,-0.046875,-0.0703125,-0.0234375,0.0625,0.0703125,-0.0390625,0.015625,-0.0546875,-0.0390625,-0.046875,-0.015625,-0.0390625,0.0234375,0.0390625,0.0625,-0.046875,-0.015625,-0.015625,0.046875,0.0546875,0.015625,-0.046875,0.015625,0.03125,0.046875,-0.0,0.0546875,0.0546875,-0.0078125,-0.0234375,-0.0078125,0.0078125,0.0,-0.0390625,-0.03125,-0.0546875,-0.0234375,0.015625,-0.0,0.0078125,0.03125,0.0859375,-0.0,-0.0234375,-0.0625,0.0078125,0.015625,-0.0234375,-0.1015625,-0.0390625,-0.03125,0.078125,-0.0234375,0.0703125,-0.0078125,-0.0625,-0.0546875,-0.0078125,0.0859375,-0.0234375,-0.03125,0.078125,0.0390625,0.0234375,-0.03125,-0.0234375,0.0390625,-0.0234375,-0.0390625,-0.046875,-0.0390625,-0.0234375,-0.0546875,0.015625,-0.0390625,-0.03125,-0.046875,-0.046875,0.0234375,-0.03125,-0.0078125,-0.0078125,-0.0390625,0.046875,0.0,0.015625,-0.0,0.0859375,-0.0546875,-0.046875,-0.0078125,0.015625,0.0078125,-0.0625,0.0078125,0.0390625,0.0703125,-0.015625,-0.015625,0.0703125,0.0,0.015625,-0.0390625,-0.0625,-0.0,-0.0078125,0.0,-0.046875,0.03125,-0.03125,0.03125,-0.015625,-0.0546875,-0.015625,0.0390625,-0.0546875,0.109375,0.046875,-0.0,-0.0703125,0.0,-0.0234375,-0.03125,0.0390625,0.03125,0.0234375,-0.0234375,-0.0078125,-0.0234375,-0.0390625,-0.0234375,0.03125,-0.0390625,-0.0,-0.015625,0.015625,-0.046875,-0.0078125,-0.015625,-0.0078125,-0.015625,0.0078125,-0.0078125,-0.046875,0.03125,-0.0234375,0.0,-0.0234375,-0.0078125,0.0078125,0.0390625,-0.015625,-0.015625,-0.0390625,0.0234375,0.0234375,-0.015625,-0.0,-0.03125,-0.046875,0.015625,0.0546875,-0.015625,0.0546875,0.09375,-0.0390625,0.03125,-0.015625,0.078125,0.078125,0.03125,-0.0,-0.03125,0.0,-0.046875,0.078125,-0.046875,0.03125,0.015625,0.046875,-0.0390625,-0.078125,-0.1015625,-0.0234375,-0.1015625,-0.0703125,0.03125,0.046875,0.015625,-0.0078125,0.0546875,-0.015625,-0.0703125,0.0234375,0.03125,0.046875,0.0234375,-0.03125,0.046875,-0.03125,0.0,-0.0,0.015625,-0.0234375,0.0546875,0.0234375,0.015625,-0.046875,0.0078125,0.0234375,0.0625,-0.0390625,-0.0078125,-0.0390625,0.0546875,-0.0703125,0.0546875,0.046875,0.015625,-0.078125,-0.03125,-0.015625,0.0703125,-0.0390625,0.0078125,0.03125,0.0,-0.0546875,-0.0390625,0.03125,-0.0234375,-0.015625,-0.0,-0.015625,-0.0390625,0.0546875,0.0,-0.03125,-0.0546875,0.046875,0.015625,0.0,0.0390625,-0.0,0.0078125,0.0234375,0.03125,0.015625,-0.03125,-0.015625,0.0390625,0.0078125,-0.0390625,-0.015625,-0.046875,-0.03125,-0.0625,-0.0390625,-0.0234375,-0.015625,-0.03125,-0.0078125,-0.0234375,0.0,-0.03125,-0.0390625,0.109375,-0.0234375,-0.0234375,-0.0390625,0.0234375,-0.03125,0.0234375,0.03125,0.0625,0.03125,-0.03125,-0.015625,0.03125,-0.046875,-0.0390625,0.03125,-0.0546875,-0.046875,-0.046875,-0.0234375,0.0625,-0.015625,0.03125,-0.015625,-0.015625,-0.0078125,-0.0,0.0,0.0234375,0.015625,-0.0390625,-0.015625,-0.0390625,0.0078125,-0.015625,-0.03125,-0.0546875,-0.015625,-0.0078125,0.03125,0.015625,-0.0078125,-0.0234375,-0.015625,0.0390625,0.09375,-0.0078125,0.03125,0.0234375,-0.0234375,-0.0078125,-0.0390625,0.015625,0.03125,0.0390625,0.0546875,-0.0390625,0.0703125,-0.0625,0.0,-0.015625,0.0234375,-0.0,0.0,0.0859375,-0.0078125,0.015625,-0.0234375,0.0078125,0.0390625,-0.0546875,0.0078125,0.0078125,-0.015625,-0.0,-0.0625,0.0078125,-0.0390625,-0.046875,-0.0703125,-0.0234375,-0.0625,0.046875,0.0390625,0.046875,-0.0703125,-0.015625,-0.0078125,0.0234375,0.0,-0.046875,-0.03125,-0.0078125,0.0625,-0.0,-0.0703125,-0.03125,0.09375,0.015625,-0.0390625,0.0234375,-0.0546875,-0.0,-0.015625,-0.0078125,-0.03125,-0.0390625,-0.0,0.0,-0.0546875,-0.0390625,0.046875,-0.0234375,-0.0390625,-0.03125,-0.03125,0.015625,0.0703125,0.015625,0.015625,0.0234375,0.015625,-0.0234375,-0.046875,-0.03125,-0.0,-0.0234375,-0.015625,0.0234375,0.0390625,-0.015625,0.0078125,0.015625,0.0,0.0078125,-0.0234375,-0.0234375,-0.0390625,0.03125,-0.0078125,-0.0,0.0390625,-0.046875,-0.03125,0.03125,0.0234375,-0.0546875,-0.03125,0.0078125,0.0390625,-0.015625,0.046875,0.0,-0.0390625,0.03125,0.046875,-0.0234375,0.015625,0.0546875,-0.0078125,-0.0,0.0078125,-0.0390625,-0.0234375,-0.0078125,-0.0390625,-0.0625,0.0390625,0.0390625,-0.015625,0.0,0.0,0.0703125,-0.046875,0.0234375,0.0625,0.0390625,0.0078125,-0.0703125,-0.0234375,-0.015625,0.0078125,-0.0234375,-0.0390625,0.0390625,-0.0546875,-0.03125,-0.0234375,-0.0234375,-0.0,-0.0234375,-0.0078125,0.0234375,0.078125,0.0234375,-0.0078125,0.03125,-0.015625,0.015625,0.0078125,-0.0234375,-0.0546875,-0.0546875,-0.0390625,-0.046875,-0.09375,0.0390625,0.0703125,0.015625,0.03125,-0.0703125,0.0625,-0.0234375,0.0703125,0.0078125,-0.0546875,-0.015625,-0.0625,-0.015625,0.1015625,0.015625,-0.0,0.03125,0.0390625,0.0,0.09375,-0.0625,-0.015625,-0.0625,0.0234375,-0.1015625,0.0,-0.0234375,-0.0546875,-0.03125,-0.0546875,-0.0546875,-0.0859375,-0.0234375,0.125,0.0859375,-0.0625,-0.015625,0.03125,-0.046875,0.046875,-0.015625,-0.015625,0.0,0.0078125,-0.0234375,0.046875,-0.03125,-0.046875,0.0,-0.0,0.0234375,0.0078125,-0.0078125,-0.0234375,0.03125,-0.0234375,0.0390625,-0.0390625,0.0,-0.0,-0.046875,0.0,-0.046875,0.0234375,-0.0546875,0.03125,-0.0546875,0.0546875,0.03125,0.078125,-0.0234375,0.0703125,-0.0546875,0.015625,-0.0234375,0.0234375,0.0234375,0.0625,0.0234375,-0.0390625,0.0078125,-0.0625,0.0078125,-0.03125,0.015625,-0.03125,-0.0234375,-0.046875,-0.015625,0.015625,-0.0625,0.0390625,-0.0234375,0.046875,-0.0546875,0.0546875,0.03125,0.046875,-0.015625,0.0390625,-0.046875,0.046875,-0.0703125,0.03125,0.0078125,0.015625,-0.0234375,0.0234375,0.046875,0.0078125,-0.015625,-0.046875,0.0546875,0.0859375,0.0390625,-0.078125,0.0546875,0.015625,0.0546875,-0.03125,-0.0,-0.0234375,0.0,-0.0625,-0.0078125,0.0625,0.078125,-0.0625,-0.03125,0.1640625,0.09375,-0.0390625,-0.0234375,-0.015625,-0.0859375,-0.03125,-0.0625,0.078125,0.015625,-0.046875,-0.0390625,-0.0234375,-0.0078125,-0.0234375,-0.0234375,0.015625,-0.03125,0.0234375,-0.0,-0.015625,0.0078125,0.015625,-0.0078125,-0.0078125,-0.03125,-0.03125,0.0,-0.03125,0.0078125,-0.0390625,0.0234375,0.0234375,0.0,-0.0078125,-0.0234375,-0.0078125,0.0078125,0.0078125,-0.0234375,-0.0703125,-0.015625,0.09375,0.109375,-0.03125,-0.015625,-0.0,-0.046875,-0.1328125,0.0625,-0.046875,-0.015625,-0.078125,-0.015625,-0.1484375,0.0234375,0.046875,0.078125,0.0078125,0.015625,-0.046875,0.1875,0.0625,-0.0390625,0.015625,-0.09375,-0.0390625,-0.0234375,0.0234375,0.03125,0.0546875,0.0234375,-0.046875,0.0078125,0.0625,-0.015625,-0.0,0.0234375,-0.0078125,0.0234375,-0.0390625,-0.046875,0.0,0.046875,0.0390625,-0.0078125,-0.03125,-0.046875,-0.03125,-0.0234375,0.0078125,-0.046875,-0.0390625,-0.0546875,0.0,0.0078125,0.015625,0.0390625,-0.0234375,0.046875,0.0,-0.015625,0.0234375,0.078125,-0.0390625,-0.0390625,-0.0625,0.078125,0.0625,0.03125,0.0078125,0.0546875,-0.0703125,-0.03125,-0.046875,0.0234375,0.0078125,-0.0078125,-0.03125,-0.0234375,-0.0078125,0.0546875,0.046875,-0.015625,0.0625,0.0078125,0.0234375,0.0234375,-0.03125,-0.0,0.078125,-0.140625,-0.0546875,0.046875,-0.0234375,-0.0,0.0546875,-0.0234375,0.03125,0.015625,-0.0625,0.03125,0.0234375,-0.046875,0.09375,0.109375,0.015625,-0.0390625,0.03125,-0.03125,0.0703125,-0.015625,-0.0078125,-0.0234375,-0.0,-0.03125,-0.0234375,-0.0078125,0.015625,-0.046875,-0.0703125,-0.0,-0.046875,0.0234375,0.015625,0.0234375,0.0390625,-0.0546875,-0.0078125,0.03125,0.0078125,0.0625,0.0234375,0.0234375,-0.0703125,-0.0390625,-0.0,-0.0390625,-0.0234375,0.0078125,-0.0390625,0.0078125,0.0234375,0.015625,-0.015625,-0.03125,-0.015625,0.03125,-0.1015625,-0.046875,0.046875,0.1484375,0.015625,-0.03125,-0.0234375,-0.0625,-0.015625,0.0234375,-0.0546875,-0.0078125,-0.03125,0.03125,-0.0390625,0.0234375,-0.015625,-0.015625,0.109375,0.015625,0.078125,-0.015625,0.0234375,0.03125,-0.0234375,-0.015625,0.0390625,-0.0078125,-0.0078125,0.0234375,0.0078125,0.0234375,-0.0703125,-0.015625,-0.0625,-0.0703125,0.0078125,-0.0078125,-0.0,-0.0390625,-0.0390625,-0.0078125,-0.0546875,-0.0390625,-0.046875,0.0234375,-0.015625,-0.0390625,-0.0234375,-0.03125,-0.0625,0.0703125,0.078125,0.0,0.015625,-0.0234375,0.0234375,0.03125,-0.0234375,0.03125,0.015625,0.0078125,0.03125,-0.0078125,-0.0859375,-0.03125,-0.015625,0.03125,-0.0546875,0.03125,0.0,0.0,-0.0625,-0.046875,0.03125,-0.0078125,0.0390625,-0.0234375,0.0234375,0.0390625,-0.0390625,-0.0078125,0.0078125,0.0234375,-0.03125,0.0,0.0078125,0.0546875,0.0,0.03125,0.0625,-0.0625,-0.0234375,-0.0546875,-0.03125,-0.0078125,-0.0546875,-0.0078125,-0.0078125,-0.0546875,-0.0390625,0.09375,0.0546875,0.078125,-0.0390625,0.1328125,-0.0625,0.0703125,0.0703125,0.015625,-0.0234375,-0.015625,-0.0390625,0.0234375,-0.0390625,0.03125,-0.0390625,0.03125,-0.0546875,0.015625,-0.0,-0.0625,0.078125,0.015625,-0.0234375,-0.03125,-0.0625,-0.046875,0.0234375,0.0234375,0.0625,-0.0234375,-0.0078125,0.015625,-0.0234375,-0.0390625,-0.046875,-0.09375,-0.0625,-0.0625,0.0703125,-0.015625,-0.0078125,-0.0703125,-0.046875,0.046875,0.046875,0.0390625,-0.0390625,0.015625,0.0078125,-0.0078125,0.0078125,0.046875,-0.015625,-0.0390625,-0.0078125,0.078125,-0.0703125,-0.046875,-0.0703125,-0.0078125,-0.0078125,0.0625,0.015625,-0.015625,-0.03125,-0.0078125,-0.015625,0.0078125,-0.0859375,0.1171875,-0.03125,-0.015625,0.0078125,-0.0625,0.0546875,0.0234375,-0.0078125,0.0546875,0.0390625,-0.0,-0.046875,-0.03125,0.0078125,0.0,0.0390625,0.0625,-0.0078125,0.0078125,-0.0,0.109375,-0.015625,0.0078125,0.0390625,0.046875,-0.0234375,-0.0703125,-0.0703125,-0.0859375,-0.015625,-0.046875,0.0234375,-0.03125,-0.0625,-0.0390625,0.03125,-0.0234375,0.046875,0.0,0.09375,-0.0234375,-0.0390625,-0.0234375,-0.03125,0.0859375,-0.046875,-0.046875,0.0390625,0.0625,-0.0234375,0.046875,-0.0546875,-0.0546875,0.03125,0.0234375,-0.0390625,-0.0390625,-0.03125,-0.0234375,-0.03125,0.03125,-0.0234375,-0.046875,0.0,-0.078125,0.0078125,-0.015625,-0.0078125,0.0,-0.03125,-0.0078125,-0.0078125,-0.0234375,-0.046875,-0.0390625,0.0,-0.03125,0.015625,0.015625,0.0390625,0.046875,-0.0078125,0.0,0.046875,0.046875,-0.0390625,-0.0078125,-0.0234375,0.0390625,0.015625,0.0078125,0.0234375,-0.03125,-0.03125,0.0078125,0.0234375,0.0078125,-0.015625,0.0234375,0.015625,-0.0703125,0.0390625,-0.0234375,-0.0390625,-0.0390625,0.109375,0.0,-0.0,-0.015625,0.0234375,-0.0,0.03125,0.0703125,-0.015625,0.0,-0.03125,0.03125,-0.03125,-0.0703125,0.0078125,0.0078125,-0.015625,0.046875,-0.0859375,0.03125,-0.0078125,-0.0390625,-0.015625,-0.0078125,0.015625,0.015625,-0.0234375,-0.0546875,-0.0,-0.0,-0.046875,-0.046875,-0.0546875,0.0390625,-0.0546875,-0.015625,0.0234375,0.046875,0.0078125,-0.015625,0.0234375,-0.0234375,0.078125,0.0390625,-0.046875,0.0546875,-0.0,0.0078125,-0.03125,-0.0390625,0.046875,0.0234375,0.0078125,0.0234375,-0.0390625,0.0234375,-0.015625,0.03125,-0.0234375,-0.03125,0.0546875,0.0234375,-0.0078125,0.0234375,0.0390625,0.03125,0.0078125,-0.046875,-0.015625,-0.03125,-0.0234375,-0.046875,0.03125,0.0,-0.0078125,0.0234375,-0.03125,-0.0,-0.015625,-0.015625,-0.0,0.046875,-0.0234375,0.0625,-0.0234375,0.0703125,0.015625,0.015625,0.0234375,0.015625,0.015625,-0.046875,-0.046875,0.0078125,0.015625,-0.0625,-0.046875,-0.0,-0.046875,0.015625,-0.0390625,-0.03125,0.0390625,0.0625,-0.015625,0.0234375,-0.0625,-0.0390625,-0.015625,0.015625,-0.03125,-0.0703125,-0.015625,-0.0078125,0.0625,0.0390625,0.0859375,-0.0234375,0.0078125,-0.046875,0.0234375,-0.015625,-0.0,-0.0078125,0.0078125,-0.03125,-0.0234375,-0.03125,0.0234375,0.03125,-0.0234375,-0.03125,0.0078125,0.0625,0.03125,0.015625,-0.0390625,-0.03125,-0.0234375,-0.015625,-0.015625,-0.0234375,0.0,-0.0078125,0.0078125,-0.0078125,0.015625,0.0234375,0.0078125,0.03125,0.015625,-0.015625,0.0234375,0.0078125,-0.0234375,-0.03125,0.0859375,0.0390625,0.0625,-0.03125,-0.0078125,0.0078125,-0.0390625,-0.015625,-0.015625,-0.0546875,-0.03125,0.03125,-0.015625,-0.0390625,0.015625,-0.015625,0.046875,-0.0234375,-0.03125,-0.015625,-0.015625,-0.0234375,-0.015625,-0.0078125,0.0234375,-0.046875,-0.0,-0.0078125,-0.0,0.015625,-0.0625,-0.0390625,0.0234375,-0.0390625,0.03125,-0.0234375,0.0390625,0.015625,0.0234375,-0.046875,-0.046875,-0.0234375,0.0078125,0.0859375,0.03125,-0.015625,-0.03125,-0.0234375,0.0078125,0.046875,0.0078125,-0.046875,0.03125,-0.046875,-0.0078125,0.078125,0.0078125,-0.0390625,-0.0234375,0.03125,-0.0078125,-0.015625,-0.0234375,-0.03125,-0.0234375,-0.0078125,-0.0703125,-0.03125,-0.0390625,-0.0078125,0.09375,0.03125,0.03125,0.046875,-0.0078125,-0.046875,0.0390625,0.0078125,-0.0078125,-0.0703125,0.078125,-0.015625,-0.09375,-0.0078125,0.015625,-0.03125,0.1328125,-0.0390625,0.0859375,0.1015625,0.0078125,0.0078125,-0.0390625,-0.015625,-0.0859375,0.078125,-0.03125,0.0390625,0.0546875,-0.015625,0.078125,0.03125,0.03125,0.0078125,-0.0390625,-0.0,-0.015625,-0.0390625,0.03125,0.015625,0.03125,-0.0234375,-0.0,0.0078125,-0.0390625,-0.078125,-0.015625,-0.0,-0.0078125,-0.0,0.0234375,0.03125,0.0078125,-0.015625,-0.0,0.0234375,-0.0,-0.046875,0.0546875,-0.015625,-0.0234375,0.0546875,0.03125,-0.0390625,-0.0234375,-0.015625,-0.0234375,-0.0546875,0.03125,0.0234375,-0.03125,0.0234375,-0.0234375,0.015625,0.0,-0.0390625,-0.0078125,-0.03125,-0.015625,0.046875,-0.0546875,0.0234375,-0.0078125,-0.015625,-0.046875,-0.0234375,0.03125,-0.03125,-0.0234375,-0.046875,-0.03125,0.0234375,0.0234375,-0.0234375,0.0078125,0.0078125,0.0078125,0.0078125,0.0234375,-0.0,0.015625,-0.0078125,0.0234375,0.0546875,-0.015625,-0.015625,-0.0078125,-0.046875,0.0390625,0.0390625,0.0546875,-0.0546875,-0.0546875,-0.03125,-0.015625,-0.0234375,-0.0390625,0.0859375,-0.046875,-0.015625,0.046875,-0.03125,0.015625,-0.0390625,-0.0625,0.1171875,-0.0625,-0.0,0.015625,0.1015625,0.015625,0.03125,-0.0703125,-0.0,-0.015625,-0.0234375,0.0234375,-0.0078125,-0.03125,0.0078125,-0.0625,-0.0234375,-0.1171875,0.0546875,0.015625,-0.0390625,0.1015625,0.078125,0.03125,0.125,-0.0,-0.015625,0.015625,-0.0078125,-0.0625,0.0078125,-0.015625,0.015625,-0.0390625,0.1171875,-0.0,0.0546875,0.03125,-0.0078125,-0.078125,0.046875,0.0234375,0.0234375,-0.0859375,-0.046875,-0.0078125,0.0703125,-0.078125,0.046875,0.0390625,-0.0078125,-0.09375,-0.0234375,0.015625,-0.0859375,-0.0546875,0.078125,-0.0,0.0390625,-0.0,-0.03125,-0.03125,-0.03125,-0.046875,0.0625,0.0078125,-0.015625,-0.078125,-0.0234375,-0.0078125,-0.0078125,0.078125,-0.1171875,0.0078125,0.0078125,0.0625,0.109375,-0.0546875,-0.0625,-0.0546875,-0.015625,0.0703125,-0.03125,-0.046875,0.015625,0.046875,-0.046875,0.015625,-0.0390625,0.03125,-0.0234375,-0.046875,0.015625,0.0703125,-0.03125,-0.03125,0.03125,0.015625,0.0078125,0.0703125,-0.046875,-0.03125,-0.0,0.015625,0.0,0.015625,-0.015625,-0.0625,0.0,-0.0078125,-0.078125,-0.046875,-0.0546875,0.0859375,0.0703125,-0.1015625,-0.0546875,0.0625,-0.0546875,0.015625,-0.0234375,-0.0234375,0.0390625,0.015625,0.0234375,-0.0234375,-0.015625,0.0859375,-0.015625,0.0234375,-0.046875,0.0234375,0.03125,-0.0,-0.0078125,-0.046875,0.0078125,-0.03125,0.0390625,0.0078125,0.0390625,-0.0,-0.046875,-0.015625,0.0078125,-0.015625,-0.0390625,-0.0234375,-0.015625,-0.046875,0.0625,0.0234375,-0.03125,-0.0,0.03125,0.0078125,0.0078125,0.046875,0.0078125,-0.0078125,-0.03125,0.015625,0.1015625,-0.0390625,-0.015625,0.015625,-0.0234375,-0.015625,-0.0078125,0.015625,0.03125,0.0234375,0.0625,-0.0625,0.1171875,-0.0703125,0.0234375,-0.0234375,-0.0390625,-0.0390625,-0.09375,0.0546875,-0.0390625,0.0234375,0.0078125,-0.03125,-0.0078125,-0.046875,-0.0234375,0.0,-0.0078125,0.0,-0.03125,0.0,-0.0234375,0.015625,0.0078125,-0.0078125,-0.0078125,0.0390625,0.0390625,0.0,0.0078125,0.0234375,0.0546875,-0.015625,-0.03125,0.0234375,0.015625,-0.0390625,-0.0390625,-0.0234375,0.046875,-0.015625,-0.015625,0.0078125,-0.0234375,-0.0234375,0.015625,-0.0390625,0.0,0.0078125,-0.0078125,-0.0234375,0.0859375,-0.0234375,-0.0078125,0.0078125,0.0078125,-0.015625,0.0390625,-0.0234375,0.0234375,-0.0390625,-0.0234375,-0.046875,0.03125,-0.0546875,-0.0,-0.0625,0.0625,-0.0546875,-0.015625,0.015625,-0.0703125,0.046875,0.03125,0.0625,-0.0078125,0.046875,-0.0234375,0.0,-0.0078125,0.0390625,-0.03125,-0.046875,0.015625,0.0234375,0.0,-0.015625,0.0390625,0.0078125,0.0546875,-0.046875,-0.0390625,0.0234375,0.0625,0.0078125,0.03125,-0.0078125,-0.046875,-0.046875,-0.0546875,0.0234375,-0.0078125,0.0703125,-0.0625,0.015625,0.0703125,-0.015625,-0.03125,0.015625,0.015625,-0.0078125,0.03125,-0.0390625,-0.015625,-0.0390625,0.109375,-0.0234375,0.046875,0.0390625,0.0234375,0.0234375,-0.0,0.015625,-0.0546875,-0.0234375,-0.0546875,-0.046875,-0.015625,-0.0703125,0.0234375,-0.0234375,-0.0234375,-0.015625,-0.03125,-0.0234375,0.0234375,0.0078125,-0.015625,0.015625,0.0234375,0.0234375,-0.03125,-0.015625,-0.03125,0.0,0.03125,-0.0390625,-0.0078125,0.0625,-0.03125,0.0234375,0.015625,-0.015625,0.0390625,0.015625,0.0234375,0.015625,0.03125,0.0078125,-0.0078125,-0.03125,0.0546875,0.046875,-0.0234375,-0.046875,-0.0078125,0.0078125,-0.015625,-0.0546875,0.0078125,-0.03125,-0.0078125,0.0234375,-0.0390625,0.046875,-0.0078125,-0.0546875,-0.0078125,-0.0390625,0.1015625,0.0390625,0.0390625,-0.0234375,-0.03125,0.0,-0.015625,0.0703125,0.0390625,-0.015625,-0.046875,-0.0,-0.0625,-0.0546875,-0.0390625,0.0234375,-0.0859375,-0.0234375,-0.0,-0.0546875,0.0078125,-0.0625,0.0078125,-0.078125,-0.015625,0.0078125,-0.015625,0.0078125,0.078125,-0.03125,0.03125,-0.0546875,-0.0390625,-0.078125,-0.0390625,-0.03125,-0.015625,0.0078125,-0.0078125,-0.0625,-0.0390625,-0.0234375,0.015625,-0.015625,-0.046875,-0.0390625,0.078125,0.1640625,0.0078125,-0.046875,-0.0,-0.0234375,-0.0078125,-0.0703125,0.0234375,0.0390625,0.03125,0.1328125,-0.0078125,-0.0078125,-0.0625,-0.015625,0.03125,0.0078125,0.0390625,-0.0390625,-0.0234375,-0.046875,-0.0078125,0.0078125,-0.015625,-0.03125,-0.0625,0.0390625,0.0234375,-0.0703125,-0.015625,-0.0078125,0.078125,-0.0234375,0.0078125,0.1015625,-0.046875,0.0078125,0.0859375,-0.046875,-0.0625,0.0078125,0.1484375,0.046875,-0.0390625,-0.078125,-0.0546875,0.0234375,0.0234375,-0.046875,-0.046875,0.0546875,-0.0,0.0546875,-0.0234375,0.03125,-0.0234375,0.0859375,0.03125,0.046875,-0.046875,-0.0546875,-0.0859375,0.0234375,0.0859375,0.1484375,-0.0625,0.0078125,0.015625,-0.0390625,-0.03125,-0.1015625,-0.09375,-0.078125,0.0,0.0078125,-0.0,-0.0546875,-0.0234375,-0.0078125,0.0234375,-0.0390625,0.0234375,-0.0703125,-0.046875,-0.046875,0.0234375,-0.015625,-0.015625,-0.0546875,-0.0078125,0.0390625,-0.03125,0.0625,-0.0625,0.0625,-0.0234375,-0.0625,0.078125,-0.078125,-0.0625,0.0,0.0390625,-0.0,0.0078125,-0.0625,0.0390625,0.0234375,-0.0078125,-0.0546875,-0.0390625,0.03125,-0.0078125,-0.015625,-0.0078125,-0.03125,0.0,0.0703125,-0.03125,0.0078125,-0.0078125,-0.0234375,-0.03125,0.0078125,0.0,0.0078125,0.0078125,-0.0234375,0.046875,-0.015625,-0.0859375,-0.0234375,-0.0390625,-0.0078125,-0.0,0.0390625,0.0859375,-0.0078125,-0.015625,0.0390625,0.0234375,0.0234375,0.0078125,-0.03125,0.0078125,-0.0390625,0.0,-0.046875,0.0234375,-0.015625,0.046875,-0.0234375,-0.03125,-0.0,0.0078125,-0.0,0.0,0.03125,0.0625,-0.015625,-0.0234375,-0.03125,-0.015625,-0.0078125,-0.0390625,0.0,0.046875,0.0546875,-0.0703125,0.046875,-0.046875,-0.03125,-0.015625,-0.0078125,0.0234375,0.015625,-0.015625,0.09375,-0.03125,-0.015625,-0.0234375,0.0078125,-0.015625,0.0078125,0.015625,0.0546875,-0.0078125,0.015625,-0.0,-0.0390625,0.0625,-0.0234375,-0.015625,0.03125,-0.0078125,-0.0,-0.0546875,0.0078125,-0.0703125,-0.03125,0.0234375,-0.015625,-0.0234375,-0.0390625,0.03125,0.046875,-0.03125,-0.0390625,0.03125,0.0390625,0.0078125,0.0234375,-0.0078125,0.140625,-0.0703125,-0.015625,0.0390625,0.015625,0.015625,-0.0078125,-0.0546875,0.1171875,0.0234375,0.1171875,-0.015625,-0.0703125,-0.0625,-0.015625,0.0078125,-0.03125,-0.03125,0.015625,-0.0234375,0.0078125,0.0390625,0.0546875,0.0390625,-0.015625,0.0078125,0.0703125,-0.0390625,-0.0234375,0.0234375,-0.03125,-0.0546875,0.1015625,-0.0234375,-0.03125,-0.0078125,0.0390625,-0.0703125,0.046875,-0.0078125,-0.0703125,0.0078125,-0.0,0.015625,-0.0703125,0.015625,0.0625,-0.0078125,0.0078125,-0.0703125,0.03125,0.03125,0.03125,-0.0,0.03125,0.0078125,0.0234375,-0.0625,0.0390625,0.03125,-0.0390625,-0.0625,0.0234375,-0.0078125,-0.0546875,-0.03125,-0.0390625,-0.0078125,-0.046875,0.0859375,-0.0,-0.03125,0.0078125,0.03125,0.03125,-0.03125,0.03125,-0.0390625,0.0078125,-0.015625,0.046875,0.015625,0.0234375,-0.0,0.0546875,-0.0234375,0.03125,0.0078125,0.0078125,-0.0546875,0.015625,0.015625,0.015625,0.0546875,0.015625,-0.015625,-0.0546875,0.0,-0.03125,-0.046875,0.0546875,0.0234375,0.0,-0.03125,-0.015625,-0.0390625,-0.046875,-0.046875,0.0703125,-0.046875,0.03125,0.0234375,-0.0390625,0.0234375,-0.0625,-0.0234375,-0.0234375,-0.046875,0.078125,-0.0,0.03125,-0.0390625,0.0,-0.0390625,-0.03125,-0.0234375,-0.03125,-0.0390625,0.03125,0.0078125,-0.015625,0.0078125,-0.0,0.03125,0.03125,0.015625,-0.0234375,0.0078125,-0.0234375,-0.0,0.0234375,-0.015625,-0.03125,-0.0390625,-0.015625,0.0234375,-0.0078125,-0.03125,0.046875,-0.0390625,0.03125,-0.0390625,-0.0234375,0.0625,-0.0625,-0.0,0.046875,0.046875,0.0390625,0.0234375,-0.0546875,0.0234375,-0.0234375,-0.046875,0.0625,-0.0234375,-0.0078125,0.0390625,-0.03125,-0.03125,-0.046875,-0.0234375,-0.015625,-0.046875,-0.0234375,-0.015625,0.0078125,-0.0546875,-0.015625,0.09375,0.0625,-0.078125,-0.0234375,0.0,0.0625,0.0390625,-0.015625,-0.03125,0.0078125,-0.03125,-0.0703125,-0.046875,-0.0390625,-0.0078125,0.0078125,0.03125,-0.0234375,0.015625,-0.03125,-0.0,0.0390625,0.0,-0.015625,-0.0234375,0.0078125,0.109375,-0.03125,-0.0078125,0.0078125,-0.046875,-0.078125,0.046875,-0.0390625,0.0078125,0.015625,0.0078125,0.0546875,-0.0625,-0.0703125,-0.03125,0.03125,0.0,-0.0390625,0.0234375,-0.0078125,-0.0703125,0.0234375,0.0234375,-0.0859375,-0.0390625,0.0,0.0390625,-0.03125,-0.015625,0.1015625,-0.109375,0.078125,0.015625,0.03125,-0.0390625,-0.015625,-0.03125,0.0078125,-0.03125,0.109375,0.015625,0.015625,0.015625,0.0,-0.0078125,-0.0,0.0234375,-0.0234375,-0.03125,-0.0078125,-0.0546875,0.015625,0.015625,-0.0078125,-0.0,-0.0234375,-0.0234375,0.0390625,0.0390625,0.03125,-0.0546875,0.03125,-0.015625,0.0625,-0.0234375,-0.0625,-0.0390625,0.0234375,-0.0625,-0.0703125,0.046875,0.015625,0.0234375,0.03125,0.03125,0.015625,0.0,0.015625,-0.0078125,-0.0390625,-0.0234375,-0.0078125,0.078125,-0.0078125,-0.015625,-0.0,-0.0390625,-0.0078125,-0.015625,-0.0234375,-0.0390625,0.015625,-0.0390625,-0.0234375,0.0078125,-0.0,-0.0,-0.046875,0.03125,0.0390625,-0.0625,-0.015625,-0.0390625,-0.03125,0.0859375,-0.0234375,0.0234375,-0.0234375,-0.015625,0.0234375,-0.015625,-0.0546875,0.0625,0.015625,0.0390625,0.0,-0.015625,-0.0078125,0.0390625,-0.0234375,0.03125,-0.0234375,0.015625,0.0,0.109375,-0.015625,-0.0078125,0.0078125,0.0,-0.046875,-0.0546875,0.0078125,-0.0390625,0.03125,-0.0234375,0.03125,-0.015625,-0.015625,-0.0390625,-0.046875,-0.0234375,-0.0078125,-0.015625,0.0078125,-0.03125,0.0078125,-0.0234375,0.0234375,-0.015625,0.0078125,0.0,-0.0390625,-0.0234375,-0.03125,0.0546875,-0.0234375,0.0078125,-0.0546875,0.0390625,0.0078125,0.0234375,-0.0,0.0546875,-0.078125,0.0,-0.015625,0.046875,0.015625,0.0390625,-0.0546875,-0.0078125,0.0625,0.125,-0.0234375,-0.0390625,0.0,-0.0234375,-0.078125,-0.0546875,0.0078125,0.0078125,0.015625,0.0234375,-0.0625,-0.0859375,-0.03125,0.015625,0.0390625,-0.0234375,0.1015625,0.09375,-0.0390625,-0.03125,-0.1015625,0.09375,0.1015625,0.03125,0.09375,0.15625,0.0234375,0.0546875,0.0234375,0.0390625,-0.09375,-0.046875,0.0546875,-0.015625,-0.0703125,-0.0390625,-0.0703125,0.015625,-0.03125,0.0390625,-0.0078125,-0.0234375,-0.0390625,-0.015625,-0.0234375,-0.0390625,0.0625,0.0625,0.0,0.109375,-0.046875,-0.03125,0.0390625,-0.0859375,0.0,-0.09375,-0.015625,0.015625,0.0546875,0.0859375,-0.046875,-0.015625,-0.0078125,0.0,0.1015625,-0.0,0.0078125,0.03125,0.0234375,-0.046875,0.0078125,-0.0546875,0.0,0.015625,-0.0625,-0.0703125,-0.015625,0.0859375,-0.0390625,-0.015625,0.0078125,0.046875,0.046875,-0.078125,0.0546875,0.0625,0.0390625,0.015625,-0.0546875,-0.015625,0.0078125,-0.046875,0.0390625,0.015625,0.0,-0.0234375,0.0546875,-0.03125,0.0390625,-0.0546875,0.09375,-0.0390625,0.0546875,-0.0078125,-0.0,-0.015625,-0.0078125,-0.0234375,0.03125,0.046875,-0.0078125,-0.0,-0.09375,0.015625,0.015625,-0.0546875,0.0546875,-0.09375,-0.0,-0.03125,-0.078125,-0.0078125,-0.0234375,-0.0078125,-0.03125,0.0,-0.03125,-0.03125,-0.03125,-0.03125,-0.0390625,0.0703125,-0.046875,0.0234375,0.015625,0.03125,-0.0234375,0.0234375,0.0234375,-0.0234375,-0.0078125,0.015625,0.0546875,0.0390625,-0.0625,-0.0703125,0.015625,0.015625,-0.0234375,-0.015625,0.0078125,0.0234375,-0.0078125,-0.0546875,0.046875,0.015625,-0.0546875,0.03125,-0.0703125,-0.078125,0.046875,-0.0078125,-0.015625,-0.0859375,0.1015625,0.0859375,-0.0625,-0.015625,0.0234375,0.0625,-0.0703125,-0.0078125,0.03125,0.03125,0.015625,0.0234375,0.0078125,0.09375,-0.0625,0.125,0.0546875,-0.015625,0.0078125,-0.0625,-0.09375,0.0,-0.0234375,-0.015625,0.0546875,-0.015625,-0.0390625,-0.015625,-0.0,-0.0,0.0625,-0.0703125,0.0234375,-0.015625,0.125,-0.0234375,-0.0078125,-0.046875,0.078125,0.1484375,0.046875,-0.046875,-0.015625,0.171875,0.0546875,0.0078125,0.0546875,-0.0546875,-0.015625,0.03125,-0.0078125,-0.1015625,-0.03125,-0.0703125,-0.046875,-0.015625,-0.015625,0.0234375,-0.0078125,-0.109375,0.1015625,0.0234375,0.03125,-0.0234375,-0.03125,0.0234375,0.015625,-0.015625,0.0,-0.015625,-0.078125,-0.015625,-0.0234375,-0.015625,-0.0078125,0.0390625,0.0546875,-0.0546875,0.0625,-0.0546875,-0.0078125,-0.046875,-0.03125,-0.03125,-0.0,-0.046875,0.1171875,0.0703125,-0.0078125,-0.015625,-0.046875,0.0078125,-0.03125,0.0078125,-0.015625,-0.046875,0.078125,-0.0546875,0.0625,-0.046875,-0.046875,0.0,-0.015625,0.015625,0.0,-0.03125,-0.015625,-0.0078125,-0.03125,-0.109375,-0.0,0.0,-0.0546875,0.078125,-0.0625,0.140625,0.0234375,0.0390625,-0.0078125,0.0546875,-0.0390625,-0.0078125,-0.03125,0.078125,-0.0078125,0.015625,-0.015625,-0.0234375,-0.109375,0.0234375,-0.1015625,-0.0234375,-0.015625,-0.0234375,-0.0234375,-0.015625,0.015625,0.0234375,0.0390625,0.0546875,0.0703125,-0.0078125,0.03125,0.0234375,0.0625,0.078125,0.0703125,-0.0546875,-0.046875,0.09375,-0.0546875,-0.0625,-0.0078125,-0.0234375,-0.0078125,0.0078125,0.015625,0.0078125,-0.015625,-0.0546875,0.046875,-0.015625,-0.0390625,0.0078125,-0.0390625,0.0625,-0.0234375,-0.046875,0.03125,0.03125,-0.0390625,0.046875,0.03125,-0.03125,-0.046875,-0.0,-0.03125,-0.0078125,0.0703125,0.0234375,-0.0078125,0.0078125,0.0234375,-0.03125,-0.0,0.0234375,0.0625,-0.03125,-0.015625,-0.03125,-0.046875,-0.0078125,-0.0546875,0.0390625,0.0,0.0,0.015625,0.078125,-0.03125,0.0546875,-0.0078125,-0.0234375,-0.0390625,-0.0234375,0.0,-0.0390625,0.0078125,-0.0390625,-0.0546875,-0.046875,0.0625,0.078125,-0.015625,-0.046875,0.046875,-0.0546875,0.0078125,0.015625,0.0703125,-0.0625,0.0234375,0.015625,0.0703125,0.0390625,-0.03125,0.015625,0.0,0.0390625,0.0390625,0.0234375,-0.0546875,-0.0234375,-0.015625,0.0546875,-0.0625,-0.0078125,-0.0234375,-0.0859375,0.046875,-0.0,0.015625,-0.0234375,0.015625,0.015625,0.03125,-0.0625,0.046875,-0.0546875,0.09375,-0.03125,-0.015625,-0.0625,-0.015625,0.0,-0.0390625,0.0703125,-0.0,0.0703125,-0.03125,-0.0546875,-0.046875,-0.0546875,-0.0390625,-0.0234375,-0.0078125,0.0078125,0.03125,-0.0078125,-0.0234375,0.0390625,0.0546875,-0.015625,-0.0234375,-0.0234375,0.0390625,-0.0546875,-0.03125,-0.0625,-0.015625,0.1328125,0.015625,0.0078125,0.015625,0.0078125,0.0,0.0234375,0.1015625,0.0234375,-0.0,-0.0078125,0.0234375,0.0234375,-0.015625,0.0234375,-0.0390625,-0.0234375,0.0078125,-0.0,0.0,-0.0,-0.0078125,-0.0390625,0.0546875,-0.03125,0.03125,-0.0,-0.0390625,-0.0,0.0078125,-0.0078125,0.078125,0.03125,-0.0390625,0.0234375,-0.078125,0.0078125,0.1015625,0.0078125,-0.0546875,0.0703125,-0.0234375,-0.0390625,-0.015625,-0.0,-0.0234375,0.046875,0.0390625,0.0859375,-0.0390625,-0.015625,-0.03125,0.03125,0.0078125,-0.0078125,-0.03125,-0.046875,0.078125,0.1015625,-0.0703125,0.078125,0.0234375,-0.0078125,0.0390625,-0.03125,-0.0625,-0.03125,-0.03125,0.0390625,0.015625,-0.0,-0.015625,0.0703125,0.015625,0.0078125,0.0546875,-0.0234375,0.0,0.0078125,-0.03125,-0.015625,0.0234375,-0.03125,-0.0078125,0.0390625,-0.0546875,-0.03125,-0.0390625,0.0390625,0.046875,0.0625,-0.0234375,-0.0546875,0.015625,-0.0078125,0.0,-0.0234375,0.0234375,-0.03125,0.015625,-0.015625,-0.0390625,-0.0234375,0.015625,0.0625,-0.0234375,0.0546875,0.0,0.0078125,0.0234375,0.046875,-0.0390625,0.0546875,-0.03125,-0.0625,-0.015625,0.0546875,-0.0234375,-0.0234375,-0.0078125,0.0390625,-0.0234375,-0.03125,0.0703125,-0.0703125,-0.015625,0.03125,-0.03125,0.046875,-0.0546875,-0.03125,-0.03125,-0.0625,0.03125,-0.0390625,-0.0390625,0.0703125,0.0703125,0.0234375,0.0234375,0.0703125,-0.0,0.0546875,0.0078125,-0.0546875,0.0078125,-0.03125,-0.03125,0.015625,-0.0703125,-0.0625,-0.0546875,0.1015625,0.0234375,0.0078125,0.078125,-0.0,-0.0546875,-0.0703125,0.03125,-0.015625,0.03125,-0.0078125,0.0078125,-0.03125,0.0234375,0.03125,0.015625,0.015625,-0.046875,0.015625,0.046875,-0.03125,-0.0,0.046875,0.0,0.0,-0.0078125,0.03125,-0.0625,0.015625,0.015625,-0.09375,0.0234375,-0.046875,0.0234375,-0.0234375,-0.0390625,0.015625,-0.0078125,-0.0,0.15625,0.015625,0.0078125,-0.0390625,-0.03125,0.1171875,-0.0546875,0.0234375,0.0625,-0.03125,-0.0078125,-0.015625,0.0234375,0.0078125,-0.0078125,-0.0234375,-0.0,-0.0703125,0.03125,0.0078125,0.0546875,0.015625,-0.046875,-0.0234375,0.0625,0.0625,-0.0234375,-0.0546875,-0.0625,0.0234375,0.0625,-0.0,-0.0078125,-0.078125,-0.0390625,0.0234375,-0.0546875,-0.0546875,0.015625,0.0390625,-0.046875,-0.03125,0.125,-0.015625,-0.0703125,0.015625,-0.0625,0.1015625,-0.0703125,-0.0078125,-0.015625,-0.015625,-0.015625,-0.0625,0.0078125,-0.0078125,-0.0390625,0.1171875,0.0546875,-0.0390625,0.0390625,0.015625,-0.0390625,0.0234375,-0.015625,-0.03125,-0.0078125,-0.015625,-0.0234375,0.015625,0.0078125,-0.03125,-0.0078125,-0.0546875,-0.03125,0.03125,0.0390625,-0.03125,0.015625,0.0390625,0.078125,-0.046875,-0.015625,0.0078125,0.0546875,-0.0625,0.03125,0.0234375,-0.0390625,-0.015625,-0.0,-0.0390625,-0.0625,-0.0390625,-0.0234375,-0.03125,-0.0234375,-0.0234375,-0.1015625,0.0234375,0.03125,-0.0546875,0.0703125,0.03125,-0.03125,0.03125,-0.046875,-0.03125,-0.109375,0.0078125,-0.0703125,-0.0390625,0.015625,-0.0390625,-0.0390625,-0.0078125,-0.0078125,0.140625,-0.0625,-0.0625,-0.03125,0.0546875,0.0390625,-0.0859375,-0.0859375,0.0078125,0.015625,-0.078125,0.0234375,-0.0078125,-0.015625,0.015625,-0.0390625,0.03125,0.03125,0.03125,0.0390625,0.0078125,-0.0390625,0.0,-0.0234375,0.046875,0.015625,0.0078125,-0.0234375,-0.046875,0.0078125,0.03125,-0.0,-0.0078125,-0.03125,0.0078125,-0.03125,-0.015625,0.0,0.0078125,-0.0234375,-0.0703125,0.03125,-0.015625,0.0078125,-0.0234375,-0.015625,-0.015625,-0.03125,0.015625,-0.015625,0.0078125,-0.046875,0.015625,-0.0,-0.015625,0.03125,-0.015625,0.015625,0.0078125,-0.0,-0.0546875,0.0234375,-0.015625,0.078125,-0.0234375,0.125,0.015625,-0.0703125,-0.0625,-0.078125,0.0234375,-0.015625,-0.0078125,0.0625,0.0703125,0.0234375,0.015625,0.0390625,0.0078125,-0.0078125,0.0078125,-0.046875,0.0234375,-0.0078125,-0.0390625,-0.0078125,0.0390625,-0.0078125,-0.03125,-0.03125,-0.0,-0.015625,-0.015625,-0.0078125,-0.015625,0.0234375,-0.0078125,0.0703125,-0.0546875,0.015625,-0.0390625,-0.0,-0.0,-0.0234375,-0.0625,-0.0703125,-0.0078125,0.09375,0.03125,-0.0390625,-0.0390625,0.0546875,-0.015625,0.09375,-0.0078125,-0.0859375,-0.0234375,-0.0078125,-0.0078125,-0.0234375,0.015625,-0.015625,0.0078125,-0.0390625,0.0234375,-0.0,-0.0234375,-0.015625,0.0234375,0.0234375,0.0234375,-0.0625,0.0234375,-0.0703125,0.0,0.078125,-0.0390625,0.046875,0.109375,0.0234375,0.078125,0.0234375,0.0234375,-0.0390625,-0.015625,-0.0078125,0.0078125,0.03125,-0.0390625,0.0078125,-0.0234375,0.0078125,0.046875,-0.046875,0.0546875,-0.03125,-0.0390625,0.03125,-0.0078125,-0.0703125,-0.0234375,0.03125,0.03125,0.0,-0.0703125,-0.0234375,-0.0078125,-0.046875,0.0625,0.0078125,0.0546875,-0.0078125,-0.0078125,-0.046875,-0.0390625,0.03125,0.046875,-0.0390625,0.0234375,-0.046875,-0.015625,0.0234375,0.0234375,-0.0078125,-0.0,-0.0078125,-0.0078125,-0.0078125,0.0625,0.03125,0.0078125,-0.046875,-0.0234375,-0.03125,0.0859375,-0.0,0.0078125,0.0546875,0.03125,-0.0703125,-0.0546875,0.015625,0.0625,-0.0390625,-0.046875,-0.0,-0.0,-0.03125,0.015625,-0.03125,0.015625,-0.015625,0.0078125,-0.03125,-0.03125,0.03125,-0.0078125,-0.0078125,-0.015625,-0.046875,-0.0234375,0.03125,-0.0390625,-0.015625,-0.0078125,0.0546875,0.0234375,-0.0078125,-0.0546875,-0.0,0.03125,-0.015625,0.03125,0.046875,0.03125,0.0078125,-0.015625,-0.0078125,0.015625,-0.046875,-0.0390625,-0.0234375,-0.0078125,-0.03125,-0.015625,-0.0078125,-0.0390625,-0.015625,0.03125,0.0234375,0.0078125,-0.0390625,-0.03125,0.0234375,0.015625,0.03125,0.0,-0.015625,-0.015625,-0.0234375,-0.0078125,0.03125,0.0390625,-0.0234375,-0.0078125,0.0234375,-0.046875,0.0234375,0.0078125,0.015625,0.015625,0.015625,0.0,0.0546875,0.0078125,0.0234375,0.078125,-0.0234375,-0.0078125,0.046875,0.015625,-0.015625,-0.0234375,0.03125,0.0078125,0.0390625,-0.0234375,-0.015625,-0.03125,-0.0390625,0.0625,-0.0078125,-0.0625,-0.0078125,-0.0078125,-0.0,-0.0546875,0.015625,-0.0234375,-0.0234375,-0.015625,0.0,-0.0078125,-0.0,0.03125,-0.03125,-0.015625,0.0390625,-0.0078125,-0.03125,-0.03125,0.03125,-0.0,-0.03125,0.0390625,-0.03125,0.0859375,0.03125,-0.0390625,0.0703125,-0.03125,0.1328125,0.015625,-0.046875,-0.0390625,0.03125,-0.0234375,-0.0390625,-0.0390625,-0.0390625,-0.0390625,-0.046875,0.015625,-0.0078125,0.0078125,-0.0625,0.09375,0.0546875,-0.015625,0.0078125,-0.0234375,0.0546875,-0.046875,-0.0,-0.03125,-0.046875,-0.0390625,-0.0234375,0.0078125,0.0390625,-0.0234375,0.0390625,-0.0078125,-0.046875,-0.046875,-0.0234375,-0.0078125,0.03125,-0.0625,0.015625,-0.03125,-0.0234375,-0.0546875,-0.03125,-0.03125,0.0234375,0.015625,0.0859375,-0.046875,0.046875,-0.015625,0.0703125,0.0859375,-0.015625,-0.0234375,0.03125,-0.0078125,0.015625,-0.0,-0.03125,0.015625,0.0078125,0.0234375,-0.078125,0.046875,-0.046875,-0.0390625,0.0234375,-0.0546875,-0.03125,-0.0,0.0078125,0.0078125,0.0234375,0.0078125,0.078125,-0.0625,-0.0078125,0.0078125,-0.0234375,0.0078125,0.0390625,0.015625,-0.0234375,-0.0078125,-0.0234375,-0.015625,-0.046875,-0.015625,-0.0078125,-0.0078125,-0.015625,-0.046875,0.03125,0.0390625,0.015625,-0.015625,-0.0234375,0.0546875,0.0546875,-0.0234375,-0.03125,-0.046875,0.0625,-0.03125,-0.0234375,0.0703125,0.03125,-0.0234375];

weight_3x3 = [-0.0234375,0.03125,-0.0078125,-0.0625,-0.0703125,-0.015625,-0.0078125,0.0234375,-0.0234375,-0.0078125,-0.0078125,-0.015625,0.0,-0.0078125,-0.0078125,0.0,-0.0078125,-0.0078125,0.0546875,-0.0546875,0.0234375,-0.015625,0.0234375,0.03125,-0.046875,-0.0078125,0.03125,0.0390625,-0.046875,0.046875,-0.0078125,0.0,0.0625,-0.015625,-0.0390625,-0.0078125,-0.0,-0.0078125,0.0546875,0.015625,-0.0859375,-0.0859375,0.0,-0.046875,-0.0859375,0.0078125,0.0078125,0.0,0.0078125,-0.0078125,0.0078125,0.0078125,-0.0078125,-0.0078125,0.078125,-0.03125,0.109375,-0.0546875,-0.015625,0.0078125,-0.0078125,-0.046875,-0.0703125,-0.0625,-0.0,-0.0234375,0.0546875,0.0390625,0.046875,-0.0,-0.046875,-0.03125,0.0078125,-0.09375,0.109375,-0.0234375,-0.1328125,0.09375,0.0078125,-0.046875,-0.0390625,-0.0078125,-0.0390625,0.0078125,-0.0078125,0.0,0.0390625,-0.0078125,0.03125,0.0234375,0.046875,0.03125,0.0390625,-0.0546875,-0.1015625,0.0078125,0.0546875,0.015625,-0.0390625,-0.0078125,0.0234375,-0.0234375,0.0,0.0625,0.015625,-0.0234375,-0.03125,-0.03125,-0.015625,0.03125,-0.015625,-0.0234375,0.015625,-0.03125,-0.0078125,0.0234375,0.0078125,-0.0234375,0.046875,0.046875,0.0546875,0.0234375,-0.0390625,0.0078125,-0.0390625,-0.0078125,0.0,0.09375,0.03125,-0.0234375,0.0078125,0.03125,0.0,-0.0234375,-0.0234375,-0.015625,0.0,-0.0,0.078125,0.015625,-0.046875,-0.0078125,0.015625,0.0078125,-0.015625,0.0078125,0.0,-0.0,0.015625,0.0234375,0.0,-0.0078125,-0.015625,-0.0,0.0078125,-0.046875,-0.046875,0.0234375,0.0234375,-0.0,-0.0234375,-0.0390625,0.046875,-0.0234375,0.015625,-0.046875,-0.078125,-0.0,-0.03125,-0.046875,-0.0234375,0.046875,-0.03125,-0.015625,0.0,0.015625,0.03125,-0.046875,-0.0390625,-0.03125,0.0390625,0.0625,0.03125,-0.03125,-0.0078125,-0.015625,0.0546875,-0.0546875,-0.078125,0.0078125,-0.0,-0.03125,0.03125,0.0078125,0.0390625,-0.0078125,-0.0078125,-0.0625,-0.0234375,-0.0234375,0.0546875,-0.015625,-0.015625,0.125,-0.0234375,-0.03125,-0.03125,-0.0078125,-0.0078125,-0.046875,0.015625,-0.0625,0.078125,-0.0078125,0.0,0.0234375,0.0078125,-0.0546875,0.015625,0.0078125,-0.0390625,0.015625,0.0078125,-0.0546875,-0.0703125,-0.0859375,0.0,0.09375,-0.0390625,-0.1171875,-0.0703125,0.046875,0.0390625,0.078125,-0.046875,0.03125,-0.078125,-0.0078125,0.0078125,-0.015625,-0.015625,-0.0,-0.0546875,-0.1328125,0.109375,0.0546875,-0.0390625,-0.0078125,-0.0859375,-0.0,0.0078125,0.03125,0.046875,-0.0234375,0.1171875,0.0234375,-0.0703125,-0.078125,0.0390625,0.0078125,-0.0078125,0.03125,-0.0,0.015625,0.0625,-0.078125,-0.1015625,0.0234375,0.0625,0.03125,0.0390625,-0.0078125,0.0546875,-0.0390625,-0.0234375,0.0,0.0,0.0078125,-0.0078125,-0.015625,-0.078125,-0.0234375,0.015625,-0.046875,0.0078125,0.0078125,0.0078125,0.0,0.015625,-0.0078125,0.0078125,-0.03125,-0.0234375,0.015625,0.015625,-0.03125,-0.0546875,-0.015625,0.0078125,0.015625,-0.0078125,0.0,0.0078125,0.0078125,0.0078125,-0.0078125,-0.0390625,0.0078125,0.0390625,-0.0390625,0.0234375,-0.0703125,-0.0546875,-0.0546875,0.0,0.0078125,0.0078125,0.0078125,-0.0,-0.0390625,-0.0234375,-0.0078125,-0.015625,-0.046875,-0.0234375,0.0078125,0.0703125,0.015625,-0.0078125,0.015625,-0.0078125,-0.0078125,0.03125,0.0078125,0.0,-0.0078125,0.0078125,0.0078125,-0.015625,0.0,-0.0,-0.0078125,-0.015625,-0.0234375,0.0859375,0.015625,-0.015625,0.0703125,0.015625,-0.0625,-0.046875,0.0390625,0.140625,0.1015625,0.0625,0.0078125,0.0234375,-0.0234375,0.046875,-0.0546875,-0.0390625,-0.0078125,-0.0390625,-0.0,-0.03125,-0.0390625,0.046875,-0.0078125,0.0390625,-0.0078125,0.0234375,-0.0,-0.03125,-0.015625,-0.015625,-0.0234375,0.0,0.0234375,0.0859375,0.0859375,0.0546875,-0.015625,0.0,-0.0078125,-0.0234375,-0.0703125,-0.046875,-0.0,0.0078125,-0.015625,0.0234375,0.03125,0.0390625,0.0078125,-0.0078125,0.0078125,-0.03125,-0.046875,0.0390625,-0.0078125,0.0078125,-0.015625,0.0234375,-0.0078125,0.015625,-0.0,-0.0078125,-0.0078125,0.015625,-0.0234375,-0.0234375,0.03125,0.1015625,0.0078125,-0.0,0.0078125,0.015625,0.0546875,-0.0,0.0078125,0.0234375,-0.046875,-0.0625,0.0078125,-0.0703125,-0.015625,0.03125,-0.0234375,0.0390625,-0.0078125,-0.0078125,-0.015625,0.0078125,-0.0078125,0.0078125,0.0,0.0234375,0.0,0.0,-0.0078125,-0.0078125,-0.03125,0.0,-0.046875,-0.0546875,0.0078125,-0.015625,-0.03125,0.0078125,0.0,-0.0234375,-0.0078125,-0.046875,0.046875,-0.046875,0.0703125,0.046875,-0.015625,0.0078125,-0.0,0.046875,0.03125,0.015625,-0.0390625,-0.0703125,0.0234375,-0.0546875,0.015625,-0.046875,-0.1015625,-0.046875,0.03125,-0.015625,0.0546875,0.0703125,0.03125,0.0,0.0078125,-0.0546875,0.015625,-0.046875,0.03125,0.0546875,-0.0078125,-0.0703125,-0.0390625,-0.03125,-0.1015625,-0.015625,-0.03125,0.046875,0.0859375,-0.0,-0.046875,0.03125,-0.015625,-0.03125,-0.03125,-0.0078125,-0.0703125,-0.046875,0.0078125,-0.0078125,0.15625,-0.015625,0.0,-0.0546875,-0.0625,0.0234375,-0.0,-0.0234375,-0.0625,0.03125,-0.03125,-0.0703125,-0.015625,0.046875,0.03125,0.0078125,-0.015625,0.0234375,-0.0078125,0.015625,0.0546875,0.03125,-0.0,-0.0546875,-0.0,-0.0078125,-0.0234375,-0.0625,0.1015625,-0.09375,-0.03125,0.0078125,-0.109375,-0.1015625,0.015625,0.1484375,0.0625,-0.0390625,-0.015625,0.0859375,-0.046875,0.015625,-0.0625,0.0859375,0.0234375,-0.0234375,0.0234375,0.109375,0.0546875,-0.015625,-0.0625,-0.0,-0.0234375,0.015625,-0.0703125,-0.0390625,-0.0546875,-0.0078125,0.0078125,-0.0859375,0.015625,0.0625,-0.015625,-0.0234375,0.03125,-0.0234375,-0.03125,-0.09375,-0.03125,0.0,-0.015625,0.015625,0.015625,0.0,-0.0078125,-0.015625,0.09375,0.0078125,0.0,0.015625,0.046875,-0.0078125,-0.0,-0.0078125,-0.0,0.0078125,-0.0078125,0.0,0.0,0.015625,-0.0078125,-0.015625,-0.0078125,-0.0390625,-0.0234375,-0.046875,0.0078125,-0.0234375,0.015625,0.015625,-0.0,-0.03125,0.0234375,0.0234375,-0.0390625,-0.015625,0.0234375,0.0,0.0,0.0234375,0.0390625,-0.015625,-0.078125,-0.046875,-0.03125,0.0,0.03125,-0.0234375,0.0078125,-0.015625,-0.0,0.0,0.0,-0.0078125,0.015625,0.0,-0.0078125,0.0234375,-0.015625,-0.015625,-0.0,-0.0078125,0.0078125,-0.015625,0.0234375,-0.03125,-0.015625,-0.0390625,-0.0390625,0.0,0.03125,-0.0234375,-0.0234375,-0.0234375,-0.0,-0.0703125,-0.0,0.015625,-0.0,-0.0546875,-0.03125,0.015625,-0.0625,-0.0,0.0078125,-0.0078125,-0.0,0.0234375,0.03125,0.015625,-0.015625,0.0703125,0.015625,-0.0625,0.0078125,-0.0,0.0390625,0.0078125,-0.0078125,-0.0390625,-0.03125,-0.03125,-0.0078125,0.0234375,-0.0078125,0.0234375,-0.0234375,-0.0390625,-0.03125,-0.015625,0.0078125,0.0078125,-0.0078125,-0.0078125,-0.046875,-0.0234375,-0.0078125,-0.0,-0.015625,-0.0,-0.015625,-0.015625,-0.0078125,-0.0234375,0.015625,-0.0,0.078125,-0.0078125,-0.0234375,-0.046875,0.078125,0.0390625,-0.0234375,0.0703125,0.0390625,0.0234375,-0.015625,0.0390625,-0.03125,-0.0,-0.0390625,-0.0859375,-0.015625,-0.015625,0.046875,0.015625,0.015625,0.0078125,-0.015625,0.0078125,-0.015625,-0.015625,-0.0078125,-0.0,0.03125,0.0078125,0.0703125,-0.03125,-0.015625,0.03125,0.0078125,-0.0,-0.03125,0.046875,-0.0,0.015625,0.0,-0.0078125,0.0234375,0.0,-0.0234375,-0.03125,0.0234375,-0.015625,-0.0625,0.0546875,0.0234375,-0.0703125,-0.03125,-0.015625,0.0078125,0.0078125,-0.015625,-0.0078125,-0.03125,-0.0546875,-0.03125,-0.03125,-0.0546875,-0.0078125,0.1015625,-0.03125,0.0546875,-0.0234375,-0.0234375,-0.0,-0.0390625,0.0078125,-0.0390625,0.015625,-0.03125,-0.0234375,0.046875,-0.03125,-0.0,-0.03125,-0.046875,0.015625,0.0234375,-0.015625,-0.046875,0.0,-0.046875,0.046875,0.0234375,-0.0078125,0.0234375,-0.046875,-0.046875,-0.0,0.0078125,-0.0390625,0.046875,0.015625,-0.0234375,-0.0703125,0.0078125,-0.0078125,0.0234375,0.046875,-0.015625,0.140625,-0.0078125,-0.015625,-0.109375,-0.0234375,-0.0234375,0.015625,-0.0625,-0.015625,-0.1015625,-0.03125,-0.0390625,0.0703125,0.078125,-0.0234375,-0.046875,-0.046875,-0.0078125,-0.015625,0.0390625,0.0390625,0.0390625,-0.1484375,-0.015625,0.078125,-0.0078125,0.0234375,0.0078125,-0.046875,0.0078125,0.0078125,-0.0390625,-0.046875,-0.0703125,-0.0234375,-0.015625,0.078125,0.0,0.0234375,-0.046875,-0.0078125,-0.0234375,-0.03125,0.0,-0.046875,0.0390625,-0.0546875,-0.03125,-0.0234375,-0.015625,-0.03125,0.03125,0.0078125,-0.0234375,0.140625,-0.0078125,-0.03125,-0.0390625,-0.0234375,-0.0234375,-0.0,0.0546875,0.0234375,-0.0078125,0.0390625,0.015625,0.015625,0.1015625,-0.046875,-0.0078125,-0.0078125,-0.0078125,0.0078125,0.0234375,-0.03125,-0.015625,-0.015625,0.0078125,-0.015625,0.0234375,-0.0,0.0078125,-0.0390625,-0.0625,-0.0234375,-0.015625,-0.015625,-0.0234375,0.0859375,-0.0625,-0.0078125,-0.046875,0.0390625,-0.0078125,-0.0078125,-0.03125,0.0234375,-0.0859375,-0.0546875,-0.0546875,-0.0234375,0.0859375,-0.0703125,0.0078125,0.046875,0.0078125,-0.0078125,-0.0078125,0.0078125,0.0,-0.015625,-0.0078125,0.0,-0.015625,-0.03125,0.03125,-0.03125,0.1328125,0.1015625,-0.078125,-0.078125,-0.0546875,-0.0078125,0.0,0.1328125,-0.015625,-0.0859375,-0.125,0.0390625,0.015625,0.1171875,0.0390625,-0.015625,-0.046875,-0.0390625,-0.03125,0.0234375,0.0,0.015625,0.140625,0.0390625,-0.015625,-0.0390625,-0.015625,-0.046875,-0.03125,0.015625,0.015625,-0.0390625,-0.0234375,0.046875,0.0390625,-0.0078125,0.0390625,0.015625,0.0390625,-0.0234375,-0.0390625,-0.078125,-0.03125,0.0703125,-0.0234375,-0.03125,0.0703125,-0.0,-0.046875,0.0078125,-0.0390625,-0.015625,0.0078125,0.0859375,-0.03125,-0.015625,-0.0,-0.0234375,0.03125,0.015625,-0.0234375,-0.0,-0.0546875,0.0546875,0.015625,-0.03125,-0.03125,-0.0,-0.0390625,0.0078125,0.03125,-0.0078125,0.0078125,0.1171875,-0.03125,0.0234375,-0.078125,-0.0625,0.0703125,-0.0625,0.0390625,-0.0390625,-0.0,-0.125,0.1015625,-0.0625,0.0703125,-0.0,-0.0078125,-0.0078125,-0.015625,0.0,-0.015625,0.015625,-0.0,-0.015625,-0.0546875,0.140625,0.046875,0.0078125,0.0234375,0.015625,-0.03125,-0.046875,-0.0234375,-0.015625,0.09375,0.0546875,-0.0390625,-0.0234375,-0.0,-0.0078125,0.03125,-0.0078125,-0.046875,-0.140625,-0.09375,-0.109375,0.0234375,0.015625,0.078125,-0.0234375,-0.046875,-0.0078125,-0.078125,-0.0078125,0.0,-0.0078125,0.0703125,-0.03125,-0.0234375,-0.015625,-0.0390625,0.0703125,0.015625,-0.1015625,-0.0234375,-0.1171875,-0.0546875,-0.0703125,0.0078125,-0.0390625,0.0078125,-0.03125,-0.0078125,0.03125,0.0234375,-0.0234375,-0.0546875,0.109375,0.015625,0.0546875,-0.0078125,-0.0234375,-0.0234375,-0.0390625,-0.015625,-0.015625,-0.09375,0.0703125,-0.03125,0.015625,0.015625,0.0703125,-0.0546875,-0.015625,-0.109375,-0.125,-0.0078125,-0.1015625,-0.0625,-0.0546875,-0.078125,0.0625,0.0234375,0.0234375,-0.0078125,-0.0234375,-0.0234375,0.0859375,-0.0546875,-0.0234375,0.015625,-0.0234375,0.0546875,-0.0234375,-0.0859375,-0.0234375,-0.0078125,0.0234375,0.0859375,-0.0078125,0.0390625,-0.03125,-0.0078125,-0.0546875,-0.03125,-0.046875,0.03125,-0.0703125,0.0859375,0.0,0.0078125,-0.0703125,-0.0703125,0.125,-0.03125,0.0234375,-0.140625,0.03125,-0.0390625,-0.125,0.0625,0.0625,0.0234375,0.046875,-0.109375,-0.109375,-0.0703125,0.015625,0.03125,0.0234375,-0.109375,0.1484375,-0.046875,0.0078125,-0.078125,-0.0078125,-0.0546875,0.03125,0.046875,-0.015625,-0.015625,0.0234375,0.0078125,-0.015625,-0.0,0.0390625,0.0703125,0.015625,-0.0078125,0.0078125,-0.0078125,0.015625,-0.0078125,-0.0,-0.0078125,0.0078125,0.0078125,-0.0,0.0078125,-0.0234375,-0.0234375,-0.0078125,-0.0390625,0.0078125,-0.0390625,0.0234375,0.0,0.0234375,-0.0,-0.0,0.0078125,0.0078125,-0.0234375,-0.046875,0.0078125,0.015625,-0.0078125,-0.0078125,0.0078125,-0.015625,-0.0625,-0.0234375,-0.0546875,0.03125,0.0078125,-0.0,-0.0078125,0.0078125,-0.0,0.0078125,-0.0,-0.0,-0.0,-0.0,-0.0234375,0.0078125,0.015625,-0.0234375,-0.015625,0.0390625,-0.046875,0.0703125,-0.0078125,0.0703125,0.015625,0.015625,0.03125,-0.015625,-0.0,-0.0078125,0.015625,-0.0078125,-0.0390625,-0.0234375,-0.0,-0.0234375,-0.015625,0.015625,0.0,-0.015625,0.0078125,-0.0078125,-0.0078125,-0.0,0.0078125,0.0078125,-0.015625,-0.0390625,-0.015625,-0.0390625,-0.015625,-0.015625,-0.015625,-0.03125,0.0078125,-0.0234375,0.015625,-0.0234375,0.0078125,-0.0078125,0.0234375,0.0,-0.015625,-0.0078125,0.015625,0.0078125,-0.0078125,0.0,0.03125,0.015625,-0.0078125,-0.0234375,0.0078125,-0.0,-0.0078125,0.03125,-0.015625,0.0234375,-0.0,-0.03125,-0.0234375,-0.0,-0.0078125,0.03125,-0.0078125,-0.03125,0.015625,0.0078125,-0.0234375,0.015625,0.0234375,0.0234375,-0.015625,-0.0078125,-0.0,0.0,-0.015625,-0.0234375,0.015625,0.0,-0.03125,0.0234375,-0.0234375,0.0,0.015625,0.0,-0.015625,0.0078125,0.0,0.0,-0.0078125,-0.0078125,-0.0078125,0.0,0.0078125,0.0078125,-0.0234375,0.015625,0.0,-0.03125,0.015625,-0.03125,0.03125,-0.0,-0.0390625,-0.0078125,0.0234375,-0.0,-0.0234375,0.0,-0.0078125,0.0390625,-0.0078125,-0.015625,-0.0,-0.0234375,-0.015625,-0.0234375,-0.0234375,-0.046875,-0.0,0.0234375,-0.03125,-0.0390625,0.046875,0.0078125,-0.0078125,-0.0234375,-0.03125,0.0078125,0.0,-0.0078125,-0.0078125,-0.0234375,0.0078125,0.0,0.0,-0.015625,-0.0234375,-0.015625,0.0234375,0.0234375,-0.0234375,0.03125,0.0390625,0.0078125,-0.0234375,0.046875,0.0078125,-0.0078125,0.03125,-0.0234375,-0.0390625,0.0078125,0.0078125,-0.03125,-0.046875,-0.0390625,0.046875,0.0078125,-0.0390625,0.0546875,0.0,-0.0234375,-0.0234375,-0.0078125,-0.0234375,-0.015625,-0.0,-0.046875,-0.0078125,0.0546875,0.0078125,-0.0390625,0.0625,0.0546875,-0.0,-0.0234375,-0.0,-0.0,0.0078125,0.0078125,-0.03125,-0.046875,-0.015625,0.0390625,0.0390625,0.0078125,0.0234375,0.0625,-0.0390625,-0.015625,-0.0234375,-0.03125,-0.03125,-0.046875,-0.015625,-0.0546875,-0.0390625,-0.0234375,-0.046875,-0.015625,0.0,-0.03125,-0.015625,-0.0078125,-0.015625,-0.03125,0.046875,0.0078125,0.03125,0.0234375,-0.03125,-0.0390625,-0.015625,0.015625,0.0078125,-0.015625,-0.0625,-0.0234375,0.015625,0.015625,-0.0078125,-0.015625,-0.0078125,0.046875,0.03125,0.0078125,-0.0390625,0.0078125,-0.0234375,-0.078125,-0.0078125,-0.0234375,0.03125,-0.0,0.0234375,0.0,-0.0,0.0234375,-0.0078125,-0.015625,0.0,-0.0078125,0.0,-0.03125,0.0390625,0.0390625,0.015625,-0.046875,-0.0078125,-0.0078125,-0.0078125,0.046875,-0.0390625,0.0390625,0.0078125,-0.03125,-0.015625,-0.015625,0.03125,0.015625,-0.0390625,0.0625,-0.0390625,-0.0234375,0.0078125,0.03125,-0.0546875,-0.046875,-0.0,0.046875,-0.0,-0.0078125,0.0,0.0,-0.0078125,0.015625,-0.0078125,-0.0,0.015625,0.0,-0.0234375,0.015625,0.0546875,-0.015625,0.015625,0.0546875,-0.0546875,0.0,0.1015625,0.0390625,0.015625,-0.0546875,-0.0625,0.0390625,-0.0703125,-0.0078125,-0.0,0.0078125,-0.0390625,-0.0546875,0.203125,-0.046875,0.0390625,-0.1328125,0.0,-0.0546875,-0.0234375,0.03125,-0.0078125,-0.0546875,-0.0546875,-0.03125,0.03125,-0.0,-0.015625,0.0859375,-0.0703125,-0.0390625,-0.046875,-0.046875,-0.015625,-0.015625,-0.0234375,0.0390625,0.0,-0.03125,0.015625,0.046875,-0.0703125,0.0078125,-0.0546875,-0.0078125,0.03125,0.03125,-0.015625,0.0078125,0.0625,-0.03125,0.0078125,0.0234375,-0.0234375,-0.0234375,-0.0078125,-0.0703125,-0.0078125,0.0078125,0.046875,0.0078125,-0.0078125,0.0390625,0.0234375,0.0390625,-0.0546875,-0.0078125,-0.0546875,-0.015625,0.0078125,0.0234375,-0.0703125,0.0546875,0.0625,0.046875,-0.0078125,-0.0234375,-0.0859375,-0.0390625,-0.0234375,-0.0,-0.0703125,-0.015625,0.0,-0.0078125,-0.0,0.0078125,-0.0078125,-0.0078125,0.0078125,0.0078125,-0.0078125,-0.0078125,-0.015625,0.0078125,-0.0390625,-0.03125,0.0234375,0.0,-0.015625,-0.03125,0.0625,0.046875,-0.0859375,0.0703125,0.046875,-0.015625,-0.0390625,0.0390625,0.078125,-0.0390625,-0.03125,0.0390625,-0.0078125,0.03125,-0.0078125,-0.0390625,0.015625,0.0859375,-0.0546875,-0.0234375,-0.0390625,0.015625,0.03125,-0.0234375,-0.015625,-0.0390625,0.0078125,0.0546875,0.046875,-0.015625,-0.0546875,-0.109375,0.046875,0.078125,-0.015625,-0.0390625,0.0703125,0.0,0.046875,-0.0625,-0.015625,-0.0078125,-0.0625,0.015625,-0.0,-0.0390625,-0.046875,0.046875,-0.0625,0.0859375,0.0,0.015625,0.0625,0.0703125,-0.015625,-0.0234375,0.03125,-0.0390625,-0.0078125,0.03125,0.0,0.015625,0.015625,-0.03125,0.0,0.03125,-0.0390625,-0.0390625,-0.015625,0.015625,0.0625,-0.0234375,0.0390625,0.046875,0.0078125,-0.015625,-0.03125,0.03125,0.0703125,0.0234375,-0.015625,-0.09375,-0.046875,0.0390625,0.1171875,0.015625,0.0078125,0.0234375,0.0546875,0.0078125,0.0234375,0.0,-0.015625,0.0625,0.03125,0.0625,-0.0859375,0.078125,-0.0546875,0.046875,-0.0390625,-0.03125,0.0625,-0.0625,0.03125,0.0703125,-0.046875,0.0234375,0.046875,0.0,0.015625,-0.046875,-0.03125,0.0078125,-0.0078125,0.015625,0.0,-0.0390625,-0.0390625,-0.046875,-0.0390625,-0.1015625,-0.0625,0.0546875,0.0546875,0.0625,0.015625,0.0,0.03125,0.03125,-0.0234375,-0.0234375,-0.046875,0.046875,-0.015625,-0.0,-0.0,0.0,-0.0078125,0.0078125,-0.0,0.015625,0.0078125,-0.0234375,-0.0390625,0.0078125,-0.0234375,-0.0234375,-0.0546875,0.046875,-0.03125,-0.015625,0.0234375,-0.0078125,-0.0390625,-0.0234375,0.0078125,0.0390625,-0.0,-0.046875,-0.0546875,-0.015625,-0.046875,0.0078125,-0.0078125,-0.0078125,-0.0,-0.015625,-0.0,-0.0078125,0.0,0.015625,0.0078125,0.0078125,0.0078125,-0.0078125,-0.0,0.0078125,-0.0078125,-0.078125,0.0078125,0.0078125,0.0078125,0.0234375,-0.0234375,-0.03125,0.0234375,0.0,-0.015625,-0.03125,-0.0390625,-0.0234375,0.03125,0.0625,0.0078125,0.0703125,0.015625,0.0546875,-0.046875,-0.0546875,0.046875,0.0078125,-0.0546875,-0.015625,-0.0625,0.0390625,-0.0625,-0.0234375,-0.0390625,0.1015625,-0.015625,-0.0546875,-0.0078125,-0.015625,0.0078125,0.0078125,-0.0,-0.0,-0.0546875,-0.0234375,0.1015625,0.0078125,-0.0234375,-0.015625,-0.015625,0.0234375,0.0390625,-0.015625,0.015625,0.0390625,0.0078125,-0.0078125,-0.0234375,-0.015625,0.0,0.03125,-0.015625,-0.046875,0.0078125,0.0078125,-0.0390625,0.0390625,-0.0078125,-0.0,-0.0078125,-0.015625,-0.015625,-0.0234375,0.03125,0.0234375,0.015625,0.0390625,0.0,-0.0234375,0.015625,0.015625,-0.0,0.0,-0.0,-0.015625,-0.03125,-0.1015625,-0.03125,0.0859375,0.015625,-0.0546875,-0.0234375,-0.0078125,-0.015625,-0.0078125,0.0078125,0.015625,0.0078125,-0.0078125,-0.0078125,0.015625,0.015625,0.0,-0.0390625,0.0234375,0.0234375,0.0078125,0.0546875,-0.0078125,0.03125,-0.015625,-0.03125,-0.0078125,0.0546875,0.0234375,-0.03125,-0.0078125,0.03125,0.015625,-0.0,-0.03125,0.0859375,0.0390625,-0.03125,-0.0234375,-0.03125,-0.0546875,-0.015625,0.0234375,-0.0078125,-0.015625,0.015625,0.09375,-0.0234375,-0.078125,0.0078125,0.0390625,-0.0625,-0.0390625,-0.0546875,0.0234375,0.03125,0.0234375,-0.0625,-0.1171875,0.109375,-0.046875,-0.046875,0.0625,-0.0546875,-0.0234375,-0.015625,-0.0234375,-0.015625,0.0234375,-0.03125,-0.0078125,-0.0390625,-0.0546875,-0.0546875,-0.015625,0.0,0.078125,0.046875,0.0859375,0.0078125,0.0078125,-0.0390625,0.046875,-0.0234375,-0.0234375,0.0234375,0.0625,0.03125,-0.0625,-0.0,0.0390625,0.03125,-0.0390625,0.0234375,0.09375,0.015625,0.078125,-0.015625,-0.0078125,0.0390625,0.046875,-0.0625,-0.046875,-0.046875,-0.0078125,-0.0859375,0.09375,0.0390625,-0.0703125,-0.0390625,0.0859375,0.0234375,-0.0078125,-0.125,-0.0703125,0.015625,0.0234375,0.03125,-0.09375,-0.078125,0.078125,-0.0234375,-0.0,0.078125,-0.0078125,-0.03125,0.03125,-0.046875,-0.125,0.03125,0.125,-0.03125,0.0,0.0546875,0.015625,-0.078125,-0.078125,-0.0625,-0.078125,-0.0546875,0.015625,-0.0390625,-0.03125,0.0234375,0.0078125,0.0078125,-0.03125,-0.0078125,0.0859375,-0.0234375,-0.0625,0.046875,0.015625,0.140625,0.046875,-0.046875,-0.09375,0.0390625,0.0,-0.015625,-0.03125,-0.0,-0.0078125,-0.0,0.0234375,-0.015625,-0.0078125,-0.0078125,-0.0078125,0.0078125,0.109375,0.0703125,-0.0078125,-0.0078125,-0.0546875,0.0234375,-0.0,0.015625,-0.0234375,0.0234375,-0.03125,0.015625,-0.0390625,-0.0234375,0.0078125,0.015625,0.0703125,-0.0,0.0625,0.015625,0.0234375,-0.0078125,-0.0703125,-0.0,-0.046875,-0.0390625,-0.0,-0.015625,0.015625,-0.0078125,0.0078125,-0.0,-0.015625,-0.0,0.0078125,0.0078125,-0.0390625,0.0625,-0.09375,0.0234375,-0.0234375,0.0,0.046875,-0.0390625,-0.0078125,0.015625,-0.0078125,0.0,-0.046875,-0.140625,-0.0859375,-0.0078125,-0.015625,-0.046875,0.015625,0.0234375,0.0078125,0.0625,-0.03125,0.0078125,0.0,-0.0234375,-0.0078125,0.0234375,0.078125,0.046875,0.0390625,0.0390625,-0.0078125,-0.015625,-0.0234375,-0.0546875,-0.0390625,-0.0078125,-0.03125,-0.0390625,0.0078125,0.046875,-0.0625,-0.03125,-0.03125,0.015625,-0.0,-0.0078125,0.03125,0.0078125,-0.03125,0.0234375,0.0078125,0.0078125,-0.0234375,0.015625,0.0078125,0.0078125,-0.0234375,-0.0,0.0078125,0.0234375,0.0,0.015625,0.0390625,-0.0234375,0.0234375,0.046875,0.0078125,-0.03125,-0.015625,-0.0078125,0.03125,-0.078125,0.109375,0.09375,-0.0703125,0.0390625,-0.0078125,-0.0546875,-0.03125,0.1328125,-0.0546875,0.0,0.0234375,0.0078125,0.015625,-0.0,-0.0234375,-0.015625,0.015625,-0.0078125,0.015625,-0.0078125,0.0234375,0.0234375,-0.0,0.0,0.0078125,0.0,0.0078125,0.0078125,0.0078125,-0.0,-0.0546875,0.0,0.015625,0.0078125,-0.046875,-0.0625,0.046875,0.1171875,-0.046875,0.0390625,0.0,-0.015625,-0.046875,0.0078125,-0.0625,-0.0390625,0.09375,-0.0234375,-0.0,-0.046875,-0.03125,-0.0390625,-0.0390625,-0.078125,-0.0703125,0.140625,0.046875,0.109375,0.015625,-0.046875,0.03125,0.03125,-0.0234375,0.0390625,-0.015625,0.0078125,-0.03125,0.03125,0.03125,-0.0234375,0.0703125,0.0390625,0.0859375,-0.0234375,-0.0625,0.109375,-0.0078125,0.09375,0.03125,-0.1015625,0.1171875,-0.0234375,0.0234375,-0.0390625,-0.0390625,-0.0,0.0546875,-0.0390625,-0.0,0.0234375,-0.046875,-0.015625,0.03125,0.015625,-0.078125,-0.03125,0.0390625,-0.0234375,-0.0390625,0.0390625,-0.0234375,-0.0859375,-0.078125,0.03125,0.078125,0.0,0.015625,-0.03125,-0.0703125,-0.0,0.0625,0.0234375,-0.0390625,-0.0234375,-0.0078125,0.1171875,-0.109375,-0.0234375,-0.0390625,-0.03125,0.0,-0.015625,-0.03125,-0.03125,0.046875,-0.0234375,0.015625,-0.03125,-0.0234375,-0.0078125,-0.015625,-0.0390625,-0.0546875,0.09375,-0.0234375,0.1015625,-0.0390625,-0.0625,-0.0,0.0078125,0.0625,-0.0546875,0.078125,-0.046875,-0.0546875,-0.015625,-0.03125,-0.0,0.015625,0.0234375,-0.03125,-0.0234375,0.0390625,0.0703125,-0.0390625,-0.046875,-0.1328125,0.015625,-0.0546875,-0.0546875,-0.046875,0.0078125,0.0078125,-0.078125,0.078125,-0.015625,-0.0,-0.0703125,-0.078125,-0.0078125,-0.0,0.0,-0.0078125,-0.015625,-0.0,-0.015625,0.0390625,0.0,-0.03125,0.015625,-0.0390625,-0.0,-0.0,0.0078125,-0.078125,-0.0078125,-0.0390625,-0.0390625,0.0078125,-0.0390625,0.0078125,0.0078125,-0.0078125,0.03125,-0.0078125,-0.0,0.015625,-0.0078125,-0.0390625,-0.078125,-0.0546875,0.0078125,0.0234375,0.015625,-0.0078125,-0.015625,0.0,0.0078125,0.0078125,-0.0078125,-0.015625,0.015625,-0.0078125,-0.0078125,-0.0390625,-0.03125,-0.0859375,-0.015625,-0.03125,0.046875,0.0390625,0.046875,0.03125,0.015625,-0.015625,-0.0,0.046875,0.1484375,0.0,-0.0,-0.0546875,0.0078125,-0.0078125,-0.0390625,-0.0234375,-0.03125,0.0234375,-0.0625,0.015625,-0.0625,0.0078125,0.0078125,-0.0,-0.015625,-0.03125,0.0625,0.015625,-0.015625,-0.046875,0.0234375,-0.1171875,-0.0546875,-0.03125,-0.0234375,-0.0703125,0.0546875,0.1015625,0.0625,0.0546875,-0.03125,-0.03125,0.0234375,-0.0,0.0,-0.0,0.015625,0.0625,0.0234375,0.015625,-0.0,-0.0234375,-0.015625,0.03125,0.03125,-0.03125,-0.015625,0.0078125,0.046875,-0.015625,-0.0,-0.03125,-0.046875,-0.0,-0.0,-0.015625,-0.0390625,-0.0390625,-0.046875,0.0234375,-0.046875,-0.0703125,0.046875,0.0078125,0.0703125,-0.0625,-0.0078125,-0.03125,-0.0703125,0.0625,-0.015625,0.046875,0.015625,0.015625,-0.0078125,0.015625,-0.0078125,0.015625,-0.015625,-0.0,-0.0078125,0.0078125,-0.0078125,-0.0234375,0.0234375,-0.0390625,-0.015625,-0.03125,-0.015625,-0.0078125,0.0234375,0.0,0.0390625,0.03125,0.03125,0.0,-0.0234375,-0.0,-0.109375,-0.0078125,-0.0,-0.046875,-0.0390625,0.015625,-0.0,0.0,-0.03125,-0.0390625,-0.09375,0.015625,-0.0234375,0.046875,-0.109375,-0.03125,-0.0625,-0.0390625,0.0546875,-0.078125,0.109375,-0.0859375,0.015625,-0.0,-0.0234375,-0.109375,0.0078125,-0.03125,-0.0234375,-0.09375,0.046875,0.0625,0.03125,0.0390625,-0.0546875,0.0234375,0.015625,-0.0546875,0.0234375,-0.0625,0.03125,-0.0,-0.0390625,-0.03125,0.0078125,-0.0390625,-0.03125,0.0390625,-0.0703125,-0.0234375,-0.0234375,-0.0234375,-0.0546875,-0.0,-0.046875,0.0546875,-0.015625,-0.0078125,0.0625,-0.0390625,0.1015625,0.0078125,-0.03125,0.03125,-0.0234375,0.0703125,-0.0703125,0.0390625,0.0703125,-0.0078125,-0.03125,-0.0,0.0078125,-0.0390625,-0.046875,-0.015625,0.0078125,0.0859375,0.03125,0.0703125,0.03125,0.046875,-0.0546875,-0.1015625,-0.0390625,0.0234375,-0.078125,-0.046875,-0.0234375,-0.1171875,-0.0625,-0.015625,0.1015625,0.015625,0.0859375,-0.0546875,-0.015625,0.0078125,-0.1015625,-0.0,0.0,0.03125,0.0625,0.0703125,-0.0078125,-0.015625,0.0390625,0.0625,0.015625,-0.0546875,0.0078125,-0.015625,0.046875,-0.078125,-0.0390625,-0.0078125,0.0234375,-0.0,0.03125,0.0,-0.03125,-0.015625,-0.046875,-0.0234375,-0.0,-0.0390625,0.0859375,0.0625,0.0703125,-0.0546875,-0.0078125,-0.015625,0.0078125,0.015625,0.0234375,-0.0078125,0.0078125,0.0078125,0.0,-0.015625,0.0078125,0.0625,-0.0078125,-0.109375,0.0625,0.015625,-0.0234375,0.0625,-0.0234375,-0.0078125,0.0234375,0.0390625,-0.03125,-0.0625,-0.0,-0.015625,0.0546875,0.0390625,0.0390625,0.109375,-0.0078125,-0.015625,-0.0625,-0.0078125,0.015625,-0.0625,0.0078125,0.0078125,0.0,-0.0,0.0078125,0.015625,0.0078125,0.0,0.0078125,0.0234375,-0.0234375,0.0078125,0.0859375,-0.046875,-0.078125,0.0859375,0.046875,-0.03125,0.0078125,0.0390625,-0.0390625,0.0703125,-0.015625,0.0703125,-0.078125,-0.0625,-0.0625,0.03125,-0.0234375,-0.0234375,0.0078125,-0.1484375,-0.0078125,0.0078125,0.09375,0.03125,0.0234375,-0.03125,-0.0078125,-0.0078125,-0.0703125,0.0,-0.046875,-0.0234375,0.0703125,-0.0,-0.0078125,-0.0546875,-0.0078125,0.0,-0.015625,-0.0,0.0546875,-0.0546875,-0.0234375,-0.046875,-0.046875,-0.0390625,0.109375,0.0234375,0.03125,0.0703125,0.0390625,-0.0234375,-0.0078125,0.015625,0.046875,-0.0390625,0.0234375,-0.0234375,-0.0234375,-0.015625,0.015625,0.046875,-0.03125,0.046875,-0.015625,-0.0234375,-0.0078125,0.015625,0.078125,0.015625,0.0390625,0.09375,-0.0234375,-0.046875,-0.0703125,-0.109375,0.09375,-0.0078125,0.015625,-0.0390625,0.0625,-0.0078125,0.0625,0.0859375,-0.015625,-0.0546875,-0.0,-0.015625,-0.0078125,0.0,-0.015625,-0.0078125,-0.015625,-0.0,-0.0,-0.0078125,-0.0,0.0234375,-0.0390625,-0.015625,0.03125,-0.015625,-0.03125,-0.0234375,-0.046875,-0.0078125,-0.0234375,-0.015625,-0.0390625,0.0234375,0.0703125,-0.046875,0.0078125,0.0390625,-0.0703125,0.015625,0.0078125,-0.0078125,-0.0234375,-0.0546875,0.0234375,0.078125,0.046875,0.1015625,-0.0,0.015625,-0.0234375,-0.015625,-0.0234375,-0.0078125,0.0546875,0.0,-0.0234375,0.0078125,0.03125,-0.0390625,-0.015625,0.015625,-0.0078125,-0.0859375,-0.0390625,0.0,-0.03125,-0.03125,-0.0546875,-0.046875,-0.0390625,0.0234375,-0.015625,0.0859375,-0.0,0.0234375,-0.0234375,-0.0234375,-0.015625,-0.015625,0.046875,-0.046875,0.046875,-0.03125,-0.046875,-0.0234375,-0.03125,0.0234375,0.03125,-0.0,-0.0078125,-0.0390625,-0.03125,-0.046875,-0.015625,-0.0625,-0.09375,-0.0546875,-0.0625,0.078125,-0.0546875,-0.015625,-0.0234375,-0.0078125,0.0625,0.0,0.1015625,0.0390625,0.0859375,0.0078125,0.015625,-0.0859375,-0.03125,0.046875,-0.03125,-0.0390625,-0.0390625,0.046875,0.1015625,0.03125,0.0859375,0.0078125,-0.015625,0.0390625,-0.0703125,-0.0703125,-0.0859375,-0.0625,-0.0078125,-0.0078125,0.015625,0.03125,-0.0625,-0.0234375,0.015625,-0.0390625,0.046875,0.0234375,0.015625,-0.015625,0.0078125,0.0546875,-0.0625,-0.03125,-0.0703125,-0.046875,-0.03125,-0.0625,-0.0390625,0.046875,-0.078125,0.109375,0.046875,-0.0,-0.0,-0.015625,-0.0390625,0.0078125,0.0390625,-0.03125,-0.0234375,-0.0234375,-0.0078125,-0.0234375,0.0078125,-0.0078125,-0.0078125,0.0,-0.0078125,0.0078125,0.0078125,-0.0078125,-0.0,-0.03125,0.015625,0.046875,0.0546875,0.078125,0.0078125,0.015625,-0.03125,-0.0078125,-0.046875,-0.015625,0.03125,0.0234375,0.015625,-0.0234375,0.0078125,-0.0234375,0.0390625,-0.078125,-0.015625,-0.0625,-0.0546875,0.0625,0.0625,0.0390625,-0.0390625,0.0,0.015625,-0.0,0.0078125,0.0078125,0.0,-0.0,-0.0,-0.0078125,-0.0,0.0078125,-0.0234375,-0.0078125,-0.0390625,0.03125,0.0546875,0.015625,-0.0546875,-0.03125,-0.0390625,0.03125,-0.0546875,0.09375,0.0234375,-0.0390625,-0.03125,-0.015625,-0.0078125,0.0390625,-0.015625,-0.0234375,-0.015625,0.078125,0.0546875,-0.0078125,-0.078125,-0.046875,0.015625,0.0,-0.0078125,0.015625,0.0546875,0.0234375,0.0078125,-0.015625,0.015625,0.0078125,-0.0,0.0078125,-0.078125,-0.0234375,0.0234375,0.0078125,0.0,-0.03125,-0.0234375,-0.0078125,-0.0234375,0.0234375,-0.015625,-0.0625,0.015625,-0.015625,-0.0078125,-0.03125,-0.0078125,0.0078125,0.0625,0.0078125,0.0,-0.03125,-0.03125,0.0,0.0078125,0.0390625,0.0,0.0625,-0.0,0.0234375,-0.0234375,-0.0078125,-0.015625,-0.03125,-0.0390625,0.015625,-0.0703125,-0.0703125,0.0390625,-0.0234375,0.0078125,-0.046875,0.0078125,-0.0234375,0.0078125,-0.0,-0.0078125,0.0390625,-0.046875,-0.015625,0.0,0.0078125,-0.015625,0.0,-0.0078125,0.0,0.0078125,-0.015625,-0.0078125,-0.0078125,-0.0,0.015625,0.046875,0.0390625,0.0390625,-0.0625,0.0,-0.0078125,-0.03125,0.0,-0.0078125,-0.03125,0.0234375,-0.0078125,-0.0390625,-0.015625,-0.0078125,-0.015625,-0.03125,-0.0625,-0.0625,0.0703125,0.0234375,0.03125,0.0078125,-0.015625,-0.0078125,0.046875,0.0703125,-0.0234375,-0.03125,0.078125,-0.0234375,-0.0,-0.03125,-0.0390625,-0.03125,-0.0078125,0.0078125,0.1171875,0.109375,-0.03125,-0.0078125,-0.03125,-0.03125,0.0234375,0.015625,-0.0234375,0.0078125,0.0078125,-0.0546875,-0.0234375,0.0,-0.0234375,-0.0078125,-0.03125,-0.0078125,0.125,0.0390625,-0.0234375,0.0234375,-0.0703125,-0.0,0.0703125,0.0703125,0.0390625,-0.0234375,0.0,-0.046875,0.015625,0.015625,-0.015625,0.0703125,-0.0234375,-0.046875,0.0234375,-0.03125,-0.0,0.0,-0.015625,-0.015625,-0.0078125,0.0078125,-0.03125,0.03125,0.1015625,0.015625,-0.046875,-0.0234375,-0.0078125,-0.078125,-0.0390625,0.0234375,-0.03125,-0.0546875,0.015625,-0.0546875,0.0,0.015625,-0.0390625,-0.015625,-0.0546875,-0.0078125,0.03125,-0.0078125,-0.0390625,-0.0078125,0.015625,-0.0625,-0.0390625,0.0625,-0.0,-0.0625,-0.0234375,-0.0078125,-0.015625,-0.0078125,0.0,-0.015625,0.0,0.0703125,-0.0703125,-0.015625,-0.0703125,-0.0078125,-0.0078125,-0.0390625,0.0234375,0.0078125,0.015625,0.0,0.0390625,0.0625,0.0234375,0.03125,-0.0234375,-0.0,-0.0546875,-0.0390625,0.0390625,-0.0234375,-0.015625,0.0078125,-0.0234375,-0.0078125,0.0078125,-0.015625,0.015625,-0.0078125,-0.0078125,-0.0078125,-0.0078125,-0.0078125,-0.015625,0.0390625,-0.0859375,0.015625,0.03125,0.0078125,-0.0625,-0.0234375,0.078125,-0.0390625,-0.03125,-0.03125,0.0546875,0.0625,-0.015625,-0.03125,0.0078125,-0.0234375,-0.0234375,-0.0,-0.0078125,0.0390625,0.015625,0.03125,0.03125,-0.0234375,-0.03125,-0.0078125,0.0234375,0.0078125,-0.0078125,0.0078125,-0.0078125,0.0,0.0078125,-0.0,-0.046875,-0.03125,-0.140625,-0.0390625,-0.015625,0.0234375,0.0078125,0.0078125,0.0234375,-0.0390625,0.0234375,-0.0625,-0.0,-0.109375,-0.0703125,-0.0234375,-0.0546875,-0.0078125,-0.03125,0.0078125,0.0078125,-0.015625,0.015625,0.03125,-0.015625,-0.0390625,-0.015625,0.015625,0.0078125,0.0078125,-0.0078125,-0.0234375,0.0234375,0.0078125,-0.0,-0.015625,-0.015625,-0.046875,-0.0234375,-0.0703125,-0.03125,0.0390625,0.109375,0.0703125,-0.0,0.0,-0.0234375,-0.0390625,-0.0078125,-0.015625,-0.0,-0.0078125,0.03125,-0.0234375,0.0078125,0.0,0.015625,-0.03125,0.015625,-0.0078125,0.0,-0.03125,-0.0078125,-0.0078125,-0.0234375,0.0,-0.015625,0.1171875,0.046875,-0.0546875,-0.0703125,-0.0078125,-0.0234375,-0.0859375,-0.0078125,0.046875,-0.078125,-0.0546875,0.1171875,-0.0390625,-0.015625,-0.0546875,-0.0390625,0.03125,0.0,0.0859375,0.0078125,0.046875,0.0078125,-0.03125,-0.0,0.0078125,-0.0078125,0.015625,-0.0,-0.015625,-0.015625,0.015625,0.015625,0.0078125,0.015625,-0.0546875,-0.046875,-0.0234375,-0.0625,-0.0234375,-0.0234375,-0.03125,0.0234375,0.0078125,-0.0390625,0.015625,-0.0078125,0.0234375,0.0390625,-0.0078125,0.03125,-0.0546875,-0.0234375,-0.0234375,-0.078125,0.015625,-0.03125,-0.015625,-0.0078125,0.015625,-0.0234375,-0.015625,-0.0234375,0.046875,-0.015625,0.0625,-0.0546875,-0.0078125,0.0078125,-0.015625,-0.0078125,-0.0078125,-0.0078125,-0.0078125,0.0,0.0078125,0.0078125,-0.0234375,0.0078125,-0.0390625,0.015625,0.015625,0.0390625,0.015625,-0.0234375,0.0234375,0.0859375,-0.0,-0.03125,0.0703125,-0.0625,0.0546875,-0.0703125,-0.03125,0.015625,0.0625,-0.0,-0.015625,-0.0078125,-0.0078125,-0.0390625,-0.0390625,0.0234375,0.0703125,-0.015625,-0.0546875,-0.046875,-0.0,0.0625,0.0078125,0.0625,0.0546875,-0.0390625,0.0078125,-0.0078125,0.046875,-0.046875,-0.0390625,0.078125,-0.0546875,-0.0625,-0.03125,-0.0078125,0.0546875,-0.0234375,0.0625,-0.0703125,-0.0390625,0.0390625,-0.0234375,-0.0703125,-0.03125,0.0078125,0.0234375,0.0,-0.078125,-0.0234375,-0.0,0.046875,0.0078125,-0.0234375,-0.0546875,-0.0234375,-0.0234375,-0.0,0.015625,0.0390625,0.0546875,0.0390625,-0.0,0.0,0.03125,-0.0,-0.03125,0.0625,-0.0234375,-0.03125,-0.015625,0.0234375,0.09375,0.0390625,0.0625,-0.015625,-0.015625,-0.0234375,0.0078125,-0.0859375,0.0,0.0078125,-0.0390625,-0.046875,-0.0390625,-0.0390625,0.0,0.0,-0.0078125,-0.03125,-0.0,0.0078125,-0.0,-0.0078125,-0.0078125,0.0078125,0.015625,0.0,-0.0,-0.0546875,0.0,0.046875,-0.0234375,-0.03125,-0.015625,0.0390625,0.015625,-0.0703125,0.03125,0.0,0.0,0.046875,0.0,-0.0546875,0.0234375,0.0234375,-0.0546875,0.0234375,0.0234375,-0.0234375,-0.0390625,0.0078125,-0.0546875,0.0625,0.015625,0.0390625,-0.015625,0.0078125,0.0,-0.0078125,0.0,-0.015625,0.0078125,0.0,-0.0078125,-0.0234375,0.0078125,-0.03125,-0.046875,0.0625,-0.0078125,-0.0234375,0.0390625,-0.0234375,-0.015625,0.046875,-0.046875,-0.0234375,-0.03125,0.0,-0.0078125,-0.0078125,0.0234375,0.0546875,-0.046875,-0.03125,0.0234375,-0.0078125,-0.046875,0.03125,-0.109375,-0.0,0.0078125,-0.0078125,-0.015625,-0.0078125,-0.0078125,-0.0078125,-0.046875,-0.0625,-0.0078125,0.046875,0.03125,0.0078125,0.0,-0.0234375,0.0546875,-0.046875,-0.0234375,0.0234375,0.0390625,0.0703125,-0.015625,-0.03125,0.015625,0.0,-0.0234375,-0.0078125,0.015625,-0.015625,0.0,-0.0234375,-0.0234375,-0.0,0.0078125,0.0078125,0.03125,-0.0078125,-0.015625,-0.0078125,0.0078125,-0.015625,0.0234375,-0.0078125,0.0078125,-0.015625,0.0078125,-0.046875,-0.0859375,0.0234375,-0.03125,-0.0078125,0.0,-0.03125,0.015625,-0.0234375,-0.0625,-0.03125,-0.0546875,0.0234375,0.0234375,-0.0234375,-0.0078125,0.0,0.0546875,0.0,-0.0234375,0.0078125,0.0078125,-0.015625,-0.015625,-0.0234375,-0.015625,0.015625,0.0,0.0078125,0.0078125,0.0,0.03125,0.0,0.03125,0.0703125,0.0,0.0703125,0.046875,-0.03125,0.0,0.03125,-0.0625,-0.046875,0.0078125,-0.0390625,-0.0078125,0.0546875,0.015625,-0.015625,-0.046875,0.03125,-0.0078125,0.0078125,-0.0390625,-0.03125,0.0546875,0.0,-0.03125,0.046875,-0.0390625,-0.0078125,0.015625,-0.0,0.0078125,0.109375,0.015625,0.0078125,0.0234375,-0.046875,-0.0078125,-0.046875,0.03125,0.03125,-0.0234375,-0.0234375,-0.015625,-0.0390625,-0.03125,0.0390625,0.015625,-0.0234375,-0.078125,0.1484375,-0.0078125,-0.0234375,-0.0234375,-0.0234375,0.015625,0.03125,0.03125,0.046875,-0.0390625,0.0234375,-0.03125,0.0078125,-0.0390625,0.03125,0.0234375,-0.0234375,-0.015625,0.046875,0.0625,-0.0859375,-0.0078125,-0.0859375,0.0390625,-0.0625,0.015625,0.015625,-0.0,-0.0234375,-0.0078125,0.0546875,0.0390625,-0.0078125,0.0078125,0.0078125,-0.046875,-0.0078125,0.046875,-0.015625,-0.1171875,-0.0234375,-0.015625,-0.0703125,0.0390625,0.046875,0.03125,0.0390625,0.046875,-0.0,-0.0234375,-0.0390625,-0.015625,0.0078125,-0.0234375,0.1015625,-0.0390625,0.015625,-0.0,0.015625,-0.0234375,-0.0078125,-0.015625,-0.03125,0.078125,-0.0625,-0.03125,0.0078125,0.0078125,0.015625,-0.03125,-0.0234375,-0.0546875,0.0703125,-0.0390625,-0.0625,-0.0234375,-0.0546875,0.0546875,-0.0546875,-0.0078125,-0.03125,0.0078125,-0.03125,0.0078125,0.0234375,-0.0390625,-0.03125,-0.0234375,0.0,-0.0078125,0.0078125,0.0,-0.0078125,0.0078125,0.0078125,-0.0078125,0.0078125,0.0078125,-0.0234375,-0.0078125,-0.0078125,0.015625,0.046875,-0.0078125,-0.0234375,-0.03125,-0.0234375,-0.046875,0.0390625,0.0625,-0.0,-0.0625,0.03125,-0.0078125,-0.0234375,-0.015625,0.0234375,-0.0234375,0.125,-0.015625,-0.1171875,-0.046875,0.0546875,0.015625,-0.015625,-0.0,0.0078125,-0.0,0.0078125,-0.0,-0.0078125,0.0,-0.0078125,0.0,-0.046875,-0.0703125,-0.0078125,-0.078125,0.03125,0.03125,-0.0234375,0.015625,-0.0234375,-0.0625,0.0234375,-0.0234375,0.1015625,-0.1171875,-0.0546875,-0.0078125,-0.015625,-0.0,-0.0234375,0.1484375,0.015625,-0.0,-0.046875,-0.0234375,0.0234375,0.015625,-0.03125,-0.0078125,0.0078125,-0.0078125,0.046875,0.046875,0.0078125,-0.046875,-0.0390625,-0.0,-0.0390625,0.046875,-0.0078125,-0.078125,-0.0234375,-0.0390625,-0.015625,0.0078125,-0.0234375,0.015625,0.0234375,0.0078125,0.0078125,0.0234375,0.0234375,0.0,0.0234375,-0.015625,0.03125,-0.015625,-0.0234375,0.0078125,0.0234375,-0.03125,-0.0078125,-0.0078125,0.015625,0.0390625,0.0,-0.015625,-0.0703125,0.015625,-0.0234375,0.015625,-0.0390625,-0.0078125,0.0390625,0.0,0.0546875,-0.0078125,-0.0078125,-0.03125,-0.0234375,-0.0078125,-0.0234375,-0.0546875,-0.0,0.046875,-0.0234375,-0.0390625,-0.03125,-0.015625,-0.0390625,-0.0,0.0078125,-0.015625,0.0078125,0.0078125,-0.0,0.0078125,-0.015625,0.0078125,0.0,-0.0,-0.015625,-0.0234375,0.0234375,0.046875,-0.015625,-0.0078125,-0.0,0.0078125,0.0625,-0.015625,-0.015625,0.0546875,0.03125,-0.0234375,-0.046875,0.0234375,-0.0078125,-0.0390625,-0.0390625,-0.0078125,-0.0234375,0.0,0.09375,-0.0234375,0.0078125,0.0,0.015625,0.015625,0.0078125,0.0234375,-0.0390625,-0.046875,-0.03125,0.0,-0.0078125,0.0234375,-0.03125,0.0859375,0.0625,0.0234375,-0.0234375,-0.0703125,-0.0625,-0.0078125,0.0234375,0.015625,-0.0703125,-0.0,0.0859375,0.015625,0.0234375,0.015625,0.0078125,-0.0,-0.0703125,-0.0703125,0.015625,0.03125,0.09375,0.046875,0.0078125,-0.0234375,-0.0390625,0.078125,-0.0703125,-0.0078125,-0.0625,0.0078125,-0.015625,0.0078125,-0.015625,0.03125,0.03125,0.0390625,-0.0078125,-0.03125,-0.015625,0.0234375,-0.0546875,-0.015625,-0.0078125,-0.0234375,-0.015625,0.0234375,0.015625,-0.0859375,-0.015625,-0.046875,-0.0,0.0703125,-0.0390625,-0.0390625,-0.0546875,0.0234375,-0.078125,0.046875,-0.03125,-0.0546875,-0.0078125,0.015625,-0.0234375,-0.0078125,-0.03125,-0.0390625,-0.015625,-0.03125,-0.015625,0.0078125,0.0,0.0234375,-0.0546875,0.03125,0.0390625,-0.0,-0.03125,-0.0234375,-0.0234375,-0.0078125,-0.046875,0.0390625,-0.0234375,0.03125,0.0078125,-0.0234375,0.015625,0.015625,0.03125,-0.0234375,0.03125,0.0546875,0.015625,-0.046875,-0.03125,-0.0234375,-0.0234375,0.0078125,-0.0234375,-0.0625,-0.0,-0.0234375,-0.0078125,-0.0234375,-0.0546875,-0.0,0.0,0.0,-0.0078125,-0.0078125,0.0,-0.0,0.0,-0.015625,-0.0234375,0.1015625,0.03125,0.0703125,0.046875,-0.0390625,0.015625,-0.015625,-0.03125,0.0078125,-0.03125,-0.0078125,0.0390625,0.0703125,-0.015625,-0.015625,-0.015625,-0.046875,0.0390625,0.1015625,0.03125,-0.0078125,-0.0390625,-0.0234375,-0.078125,0.0234375,-0.0,-0.0078125,-0.0078125,0.0,-0.0078125,0.0,0.0,0.0078125,0.0078125,0.0078125,-0.0390625,0.0546875,-0.03125,0.046875,0.0234375,-0.0390625,0.0078125,0.1015625,-0.0,-0.015625,0.03125,0.015625,-0.0859375,-0.0,-0.0234375,-0.03125,0.0078125,-0.015625,-0.0078125,0.0546875,-0.0078125,-0.0625,0.015625,-0.0078125,0.03125,0.015625,-0.015625,-0.046875,0.0,-0.0,-0.0,0.0390625,0.015625,-0.046875,-0.0390625,-0.0078125,-0.03125,-0.0234375,-0.0390625,0.0390625,-0.0078125,-0.03125,-0.0390625,-0.0390625,-0.03125,-0.0546875,-0.015625,-0.046875,-0.03125,-0.03125,-0.015625,-0.0,0.0703125,-0.0,0.0078125,0.046875,-0.015625,-0.0078125,-0.0078125,-0.0,-0.0234375,-0.0546875,0.0234375,-0.0078125,0.015625,-0.0234375,-0.015625,0.0078125,0.015625,0.0,0.0234375,0.03125,-0.0390625,-0.0546875,-0.0078125,0.0,0.015625,0.0078125,0.078125,-0.03125,-0.03125,0.015625,-0.0078125,-0.0,-0.0625,0.046875,0.0,0.015625,0.046875,0.0078125,0.0078125,-0.0078125,0.0078125,0.0,0.0,-0.0078125,-0.0,0.0,0.0,-0.0234375,-0.0,-0.0078125,-0.0,0.0234375,-0.0,0.015625,0.078125,0.0078125,0.0078125,-0.015625,0.015625,-0.0234375,-0.015625,-0.0234375,-0.0703125,-0.046875,-0.0234375,-0.0078125,-0.0234375,-0.015625,0.0234375,-0.0234375,-0.03125,0.046875,-0.015625,-0.015625,-0.0390625,-0.078125,-0.015625,0.03125,-0.0703125,-0.0078125,-0.0078125,-0.0390625,0.0,0.0546875,0.03125,-0.03125,-0.0078125,-0.015625,-0.0078125,0.0078125,-0.0234375,0.0234375,-0.0078125,-0.03125,0.0234375,0.03125,-0.0078125,-0.0546875,0.03125,0.046875,-0.0,-0.0390625,-0.03125,-0.0078125,0.03125,-0.0390625,-0.0078125,0.109375,-0.015625,-0.03125,0.0234375,-0.0234375,-0.0078125,-0.0,-0.015625,-0.015625,-0.015625,0.046875,-0.0,-0.0390625,-0.03125,-0.0078125,0.0234375,0.0390625,-0.015625,-0.0703125,0.0078125,0.046875,0.0078125,0.015625,0.03125,-0.046875,-0.0390625,-0.03125,-0.0703125,0.015625,0.0390625,-0.0390625,0.046875,-0.015625,0.0390625,-0.015625,0.0078125,-0.015625,-0.015625,0.0625,-0.0234375,-0.0390625,-0.03125,0.0625,-0.0625,-0.0390625,-0.03125,-0.0390625,-0.03125,-0.0234375,-0.0078125,-0.015625,0.0,0.0859375,-0.0234375,-0.015625,-0.0,-0.0234375,0.015625,0.0234375,0.015625,-0.0703125,0.015625,-0.0390625,0.0,-0.0078125,0.0234375,-0.0,-0.0703125,-0.015625,-0.0625,0.0078125,-0.03125,-0.03125,0.03125,-0.015625,-0.03125,-0.046875,-0.0703125,-0.0078125,-0.0234375,-0.046875,-0.0078125,0.046875,0.09375,0.0078125,0.0078125,0.0078125,-0.0078125,-0.0078125,-0.0078125,-0.0078125,0.0078125,0.015625,-0.0546875,0.046875,0.0546875,-0.03125,0.0234375,-0.046875,-0.046875,0.015625,0.0234375,-0.0078125,0.0390625,0.078125,0.0390625,0.0546875,-0.0234375,-0.0390625,-0.015625,0.0859375,-0.0546875,0.0,-0.0390625,0.03125,0.046875,-0.0546875,0.0078125,0.0625,-0.0078125,-0.0,-0.0078125,0.0078125,0.0,0.0078125,-0.0,-0.0078125,-0.015625,-0.0078125,0.0078125,-0.0859375,0.078125,-0.015625,-0.015625,-0.0625,-0.0234375,-0.046875,0.0390625,0.03125,-0.046875,-0.015625,-0.015625,-0.046875,-0.0859375,0.0,0.03125,-0.0234375,-0.0078125,-0.015625,0.0,0.0703125,0.0859375,-0.0390625,-0.0078125,-0.0078125,-0.046875,0.0,0.0390625,-0.046875,-0.0390625,0.0390625,0.015625,0.0234375,0.0234375,-0.03125,-0.0,0.0703125,0.0078125,-0.1015625,0.0078125,0.03125,-0.0,0.0546875,0.0390625,0.0,0.0078125,-0.0078125,0.0078125,0.0078125,-0.03125,-0.0234375,-0.0546875,-0.0390625,-0.0,-0.0234375,0.0390625,0.0390625,-0.0078125,-0.015625,-0.015625,0.0078125,0.0,-0.0,-0.0234375,0.0,0.0,-0.015625,0.1640625,-0.0,-0.03125,0.0078125,0.0234375,-0.0078125,-0.125,-0.0703125,0.0859375,0.078125,-0.046875,-0.09375,-0.0703125,-0.0078125,0.0234375,0.0234375,-0.03125,0.0234375,-0.0390625,-0.046875,-0.0078125,-0.046875,-0.0078125,-0.0234375,0.0078125,0.0078125,-0.03125,0.015625,-0.0078125,0.0078125,-0.0078125,-0.03125,0.015625,-0.0625,-0.015625,0.015625,-0.0234375,0.0390625,-0.0078125,0.015625,0.046875,0.0390625,-0.0,-0.0078125,0.0078125,0.0,-0.0,-0.0,0.0234375,-0.0390625,-0.0546875,-0.03125,-0.015625,0.0078125,0.0078125,-0.0390625,-0.03125,0.015625,0.0390625,-0.015625,-0.015625,0.03125,0.0,0.0703125,0.015625,0.015625,-0.0078125,-0.03125,-0.0390625,-0.0390625,-0.03125,0.0234375,-0.0,-0.046875,0.015625,0.03125,0.0078125,0.0390625,-0.09375,0.0234375,0.0,-0.046875,-0.0546875,0.015625,-0.0078125,-0.015625,-0.0390625,0.1640625,-0.0625,-0.046875,-0.09375,0.0078125,0.046875,0.0078125,-0.046875,-0.015625,0.0,-0.0,0.0390625,0.0,-0.0390625,0.0859375,-0.0546875,-0.0390625,0.0078125,-0.0625,-0.0546875,0.0625,0.015625,0.03125,0.03125,-0.0390625,-0.0234375,-0.03125,-0.0234375,0.0859375,-0.1171875,0.0234375,-0.046875,-0.0390625,0.046875,-0.0,0.0625,-0.09375,0.03125,-0.015625,0.0859375,0.078125,-0.09375,-0.0625,-0.0078125,-0.0390625,-0.0234375,-0.046875,0.0390625,0.0546875,0.078125,-0.0390625,0.0,-0.0625,0.0,0.09375,-0.078125,-0.0,-0.109375,0.1015625,-0.0625,0.0703125,0.0546875,-0.0078125,-0.0234375,0.0078125,-0.0078125,-0.0390625,0.0,0.0546875,0.0390625,-0.0703125,-0.0234375,0.046875,-0.0625,-0.0390625,-0.046875,-0.0078125,-0.0625,0.078125,0.015625,0.0703125,-0.0234375,0.0078125,-0.0078125,-0.0078125,-0.0390625,-0.046875,-0.0234375,-0.015625,-0.0,-0.015625,0.0,0.015625,-0.0,0.0078125,0.0078125,-0.0,-0.0390625,-0.0234375,-0.0625,-0.0078125,-0.078125,-0.0703125,0.03125,0.0,0.015625,0.0,-0.03125,-0.0390625,0.0078125,0.0078125,-0.0234375,-0.03125,0.0,0.0078125,0.0078125,0.0234375,-0.046875,-0.078125,0.0078125,-0.015625,-0.03125,0.015625,-0.0078125,0.0078125,0.015625,0.0078125,0.0,-0.0078125,-0.0,-0.0078125,0.0078125,-0.0078125,-0.0625,-0.0546875,-0.0703125,-0.015625,0.015625,-0.0625,-0.0234375,-0.0078125,0.015625,0.0078125,-0.015625,-0.0,-0.015625,0.0390625,0.0703125,-0.0078125,0.0234375,0.0234375,-0.03125,-0.0,0.0078125,0.0390625,0.0390625,0.0703125,0.0390625,-0.0234375,0.0078125,-0.03125,0.0078125,0.0234375,-0.0078125,-0.03125,0.0390625,0.0,0.0234375,0.0234375,0.0390625,-0.0546875,-0.015625,0.0,0.046875,0.015625,-0.0234375,-0.015625,-0.0078125,-0.0078125,0.03125,-0.0234375,-0.0234375,0.0078125,-0.0234375,-0.015625,-0.015625,0.0,-0.015625,-0.015625,0.0390625,-0.0078125,-0.0390625,0.0078125,-0.0234375,-0.0078125,0.0234375,0.0,0.0,-0.0078125,-0.03125,-0.046875,-0.0078125,-0.0234375,0.015625,-0.015625,0.03125,-0.0546875,0.03125,0.0234375,-0.0078125,0.0703125,-0.0234375,-0.0234375,-0.0546875,0.046875,-0.0234375,-0.0390625,-0.0234375,0.0234375,-0.03125,-0.03125,0.0078125,-0.0,-0.0078125,-0.0078125,0.0078125,0.0234375,-0.0,-0.0078125,-0.015625,0.0078125,-0.015625,-0.015625,0.03125,0.0390625,-0.015625,-0.015625,-0.03125,-0.0234375,-0.0078125,0.015625,-0.0390625,0.03125,0.03125,-0.0234375,0.015625,-0.0078125,0.0546875,0.0,0.0078125,-0.03125,0.0390625,0.0,-0.03125,0.015625,-0.0,-0.0078125,-0.0546875,-0.0078125,-0.0078125,0.09375,-0.03125,0.015625,0.0703125,-0.0859375,-0.046875,-0.0390625,-0.03125,-0.015625,-0.0234375,-0.0,0.0,-0.0078125,0.0,0.0,0.0390625,0.0078125,-0.0859375,0.109375,-0.0625,-0.0078125,0.0078125,-0.0546875,0.0625,-0.0234375,-0.0078125,0.125,-0.015625,0.046875,-0.0546875,-0.015625,-0.078125,-0.0546875,-0.015625,0.0,-0.015625,0.015625,0.0078125,-0.046875,-0.0,-0.0390625,-0.0078125,0.0390625,0.015625,-0.0,0.0,-0.0546875,0.0390625,0.0078125,0.0390625,0.046875,0.0625,0.0703125,-0.03125,-0.015625,0.03125,0.015625,0.0234375,0.0234375,-0.0625,-0.0546875,-0.046875,0.0625,-0.0234375,0.0390625,0.0078125,0.0234375,0.0234375,-0.046875,0.03125,-0.0234375,0.03125,0.0,0.0078125,-0.0234375,-0.0546875,-0.015625,0.0078125,0.0234375,0.0078125,0.0078125,-0.0234375,-0.0078125,-0.0,-0.0546875,0.0,0.046875,-0.046875,0.0546875,-0.046875,0.140625,-0.03125,-0.0390625,-0.0390625,-0.0390625,0.0078125,-0.03125,-0.0390625,0.1015625,0.0390625,-0.0234375,-0.046875,-0.046875,0.0546875,0.0078125,0.0234375,-0.0546875,-0.03125,-0.0546875,-0.0078125,-0.0625,0.0,-0.0078125,-0.046875,0.1015625,0.0234375,0.0078125,0.0,0.0078125,-0.0,0.0078125,0.0078125,-0.015625,0.0,-0.0078125,-0.0546875,0.046875,0.046875,-0.0625,-0.0234375,0.0390625,-0.0234375,0.0,-0.0234375,0.0078125,0.0625,0.0078125,-0.0390625,-0.03125,-0.03125,-0.0234375,-0.0234375,0.0078125,0.1015625,0.0546875,-0.046875,-0.0078125,-0.0546875,-0.0234375,0.0078125,-0.0078125,0.03125,-0.0,-0.0078125,0.0,-0.0,-0.015625,0.0078125,-0.0078125,-0.0078125,0.0078125,0.0,0.046875,0.0078125,-0.0,0.0390625,-0.046875,-0.015625,-0.03125,0.0234375,0.0390625,-0.046875,0.0546875,-0.0546875,-0.0703125,-0.0390625,-0.03125,-0.0234375,-0.0390625,0.171875,0.015625,-0.046875,-0.03125,0.015625,-0.0390625,-0.015625,-0.03125,-0.0078125,-0.0078125,0.0078125,-0.015625,-0.03125,0.0234375,0.0234375,-0.046875,-0.015625,-0.0078125,-0.0703125,0.0546875,0.015625,0.0625,0.015625,-0.0390625,-0.0546875,-0.0234375,-0.03125,0.0625,0.0,-0.0546875,-0.0,0.0390625,-0.0078125,0.015625,0.0078125,0.0,0.03125,-0.015625,-0.015625,-0.0078125,-0.015625,0.0078125,-0.015625,-0.015625,-0.0390625,-0.0,0.0234375,-0.0078125,-0.046875,-0.0078125,0.015625,0.03125,-0.015625,-0.0234375,-0.0,-0.046875,-0.0,0.015625,-0.03125,-0.046875,-0.0390625,0.0546875,-0.015625,0.046875,0.046875,-0.0625,-0.0859375,-0.046875,-0.0,0.0390625,-0.015625,0.0,0.0,-0.0078125,-0.0078125,0.0234375,-0.0,0.0078125,-0.0078125,-0.0078125,0.0234375,0.0078125,0.0078125,0.0078125,-0.0390625,0.0390625,-0.03125,-0.0234375,0.0078125,0.0,-0.0390625,0.015625,0.0625,-0.0390625,0.0234375,0.0078125,-0.0,-0.0078125,-0.015625,0.0625,-0.0,-0.0234375,0.015625,-0.046875,-0.0234375,-0.0078125,0.015625,0.015625,-0.046875,0.046875,0.0625,0.046875,-0.0234375,-0.0546875,-0.015625,-0.0234375,0.0,0.0078125,-0.0390625,0.0,-0.1015625,0.0078125,0.0078125,-0.015625,0.015625,0.0234375,-0.0234375,0.0234375,-0.0546875,0.0546875,-0.0859375,-0.0234375,0.015625,0.0078125,0.03125,0.171875,-0.0390625,0.0078125,-0.0078125,-0.0703125,-0.03125,-0.0078125,0.015625,0.015625,0.0,0.0234375,-0.0390625,0.0859375,0.0078125,-0.0625,-0.0859375,-0.015625,-0.03125,-0.0,-0.0859375,0.0,0.09375,-0.140625,0.0234375,0.0234375,0.0078125,-0.015625,-0.0078125,0.0078125,0.0625,-0.03125,-0.0,-0.0078125,-0.0234375,0.0078125,0.046875,-0.0078125,0.046875,-0.046875,-0.0234375,-0.015625,0.0546875,0.03125,-0.0,-0.0234375,0.0234375,-0.0234375,0.0859375,0.0703125,-0.046875,0.046875,-0.015625,-0.046875,-0.015625,0.046875,0.0625,0.03125,0.046875,0.0078125,-0.015625,-0.046875,-0.03125,-0.046875,-0.0078125,-0.015625,-0.0078125,0.0390625,-0.0234375,0.015625,-0.03125,-0.046875,0.0078125,-0.0546875,-0.0390625,0.0078125,-0.0078125,-0.03125,-0.0234375,0.0078125,0.0078125,0.03125,-0.046875,0.0234375,-0.0234375,-0.046875,-0.0078125,-0.03125,0.0625,0.046875,-0.0,-0.0078125,-0.015625,0.0078125,-0.0078125,-0.0078125,-0.0078125,-0.0,0.0078125,-0.0078125,0.0234375,-0.046875,-0.0625,-0.0234375,-0.0625,0.0625,0.125,0.015625,-0.046875,-0.0390625,0.0625,-0.0703125,0.0546875,-0.0546875,-0.0390625,0.0234375,0.0625,-0.015625,0.0546875,-0.03125,-0.0546875,-0.0703125,-0.03125,-0.0625,-0.0390625,-0.09375,-0.0703125,0.0,0.0078125,-0.0,-0.0,-0.0,-0.0078125,0.0078125,0.0,0.0,-0.1171875,0.0234375,-0.0546875,-0.0078125,0.0390625,-0.09375,-0.0078125,0.078125,-0.046875,-0.0390625,-0.046875,0.0390625,0.03125,-0.0625,-0.0234375,-0.03125,0.015625,-0.0078125,0.0390625,0.0,-0.015625,-0.0390625,-0.078125,-0.015625,-0.0078125,-0.03125,-0.1015625,-0.0390625,-0.0390625,0.015625,0.046875,0.015625,0.0390625,0.0,-0.0,-0.0078125,-0.0625,0.0078125,0.015625,-0.0078125,0.0546875,-0.03125,-0.0078125,-0.015625,0.015625,-0.015625,-0.0234375,0.015625,-0.0234375,-0.015625,-0.0,-0.0234375,-0.0390625,0.0078125,-0.015625,-0.0078125,0.0078125,0.0546875,-0.0234375,-0.015625,-0.0234375,-0.03125,0.0078125,0.0078125,0.0234375,-0.0,0.0078125,-0.0234375,0.0625,-0.03125,0.0390625,-0.0078125,-0.046875,-0.0390625,-0.0,0.078125,0.0859375,-0.03125,0.0078125,-0.0390625,0.0390625,-0.0625,0.0078125,0.0,-0.0234375,-0.0078125,-0.03125,0.03125,-0.0703125,0.03125,0.0,0.0,0.0234375,0.015625,0.0390625,0.0078125,-0.0,0.015625,0.0,0.0,-0.0078125,-0.0390625,0.015625,0.0078125,-0.046875,0.0390625,0.0,-0.0703125,-0.015625,0.0390625,-0.09375,-0.015625,0.046875,-0.109375,-0.078125,0.109375,-0.0234375,0.015625,-0.03125,0.015625,0.0,-0.0234375,-0.03125,-0.0234375,-0.015625,-0.0078125,0.03125,0.0546875,0.015625,0.0,0.0,0.0234375,-0.0390625,-0.0625,0.0390625,-0.125,-0.0703125,-0.0078125,0.0234375,-0.046875,-0.0546875,0.15625,0.0,-0.0625,-0.015625,-0.078125,-0.03125,-0.0625,-0.0390625,0.0625,0.0078125,0.0234375,0.015625,0.0,-0.03125,0.078125,-0.046875,-0.0390625,0.0859375,0.09375,0.1328125,0.0078125,-0.0234375,-0.0546875,-0.03125,-0.0234375,-0.0234375,0.015625,0.078125,-0.0234375,-0.015625,-0.0234375,-0.078125,-0.03125,-0.03125,0.0703125,0.0234375,0.015625,0.046875,0.046875,0.015625,0.0546875,0.0390625,-0.0234375,-0.0625,0.0078125,-0.0390625,0.0234375,0.0078125,0.109375,-0.0234375,0.0234375,0.0078125,-0.015625,0.0703125,-0.03125,-0.03125,0.0234375,0.046875,0.0,0.0078125,-0.046875,0.09375,0.0703125,-0.09375,0.0703125,0.0234375,-0.0078125,-0.0234375,0.0625,0.0703125,0.03125,0.0546875,-0.0078125,0.03125,0.015625,0.0625,0.015625,-0.015625,-0.046875,-0.1015625,0.0390625,0.03125,0.0,0.0546875,0.0078125,-0.03125,0.0234375,-0.03125,-0.03125,-0.078125,-0.0,-0.0859375,0.0078125,0.03125,0.03125,0.0078125,-0.0390625,-0.0078125,-0.0078125,0.0,-0.0390625,-0.015625,-0.0078125,-0.0078125,0.0078125,0.0078125,0.0234375,0.0078125,0.0078125,-0.0,-0.0078125,-0.03125,-0.0390625,-0.015625,-0.015625,0.015625,0.0078125,0.03125,-0.0078125,0.0078125,-0.03125,-0.015625,-0.015625,0.0078125,0.0,-0.0234375,-0.015625,-0.0390625,-0.015625,-0.0390625,-0.015625,0.0078125,0.03125,-0.0234375,-0.015625,-0.0234375,0.03125,0.0,-0.0,0.0078125,0.0078125,0.0078125,0.0078125,-0.0078125,0.0078125,-0.0078125,-0.0,0.0,0.0234375,-0.0234375,-0.0078125,0.0703125,-0.015625,-0.015625,0.0390625,0.0078125,-0.015625,-0.0546875,0.0078125,-0.0,-0.0078125,0.0078125,-0.015625,0.015625,-0.0,0.015625,-0.0625,-0.015625,0.0546875,0.03125,-0.03125,-0.03125,-0.0234375,-0.015625,-0.03125,0.0078125,0.0078125,0.03125,-0.0078125,-0.0,-0.0,-0.0234375,0.015625,-0.0234375,-0.015625,-0.015625,-0.0390625,0.0,-0.015625,-0.015625,-0.0,-0.0234375,-0.0078125,-0.03125,-0.0078125,0.0078125,-0.015625,-0.0234375,-0.0078125,-0.015625,0.0078125,0.0078125,0.0,-0.015625,0.0234375,0.0546875,0.0,-0.015625,0.015625,-0.0078125,0.03125,0.015625,-0.0078125,0.046875,-0.0,0.0078125,-0.0078125,0.0234375,0.0078125,-0.03125,0.03125,0.0,-0.015625,-0.03125,0.0,-0.0390625,-0.03125,-0.015625,0.03125,0.0625,-0.0078125,0.0,-0.03125,-0.0234375,-0.015625,-0.015625,-0.0078125,-0.0,-0.0078125,-0.0078125,0.0078125,0.0078125,-0.015625,-0.015625,0.0078125,0.0078125,-0.03125,-0.0546875,0.0078125,0.03125,0.046875,0.0078125,0.015625,-0.015625,0.0078125,-0.0703125,0.0078125,-0.0234375,-0.015625,0.03125,-0.0078125,-0.0078125,-0.015625,0.0,0.03125,0.0,-0.0234375,0.0,-0.0390625,0.015625,-0.0390625,0.03125,-0.0078125,-0.0078125,-0.0078125,-0.0,0.0234375,0.0,0.015625,-0.0,0.0078125,-0.0078125,-0.046875,0.0078125,-0.0234375,0.0703125,-0.0234375,-0.0390625,-0.0234375,0.0078125,-0.0078125,0.03125,-0.0078125,-0.0078125,-0.0390625,0.0078125,-0.0,-0.0078125,-0.0234375,-0.03125,0.0390625,-0.03125,-0.03125,0.0078125,0.0859375,0.0078125,-0.0234375,-0.0,-0.046875,-0.0859375,-0.03125,-0.0,0.0234375,0.0390625,-0.0078125,0.0390625,-0.0078125,-0.0078125,-0.0234375,-0.015625,-0.0078125,-0.046875,-0.015625,-0.015625,-0.0234375,-0.0078125,-0.0234375,0.0234375,0.015625,-0.0,0.0078125,-0.0390625,-0.0,-0.015625,-0.0234375,-0.0078125,0.046875,0.046875,0.0,0.046875,-0.015625,0.015625,-0.0390625,-0.0546875,-0.0234375,-0.03125,-0.015625,-0.015625,-0.0,0.0,0.0390625,-0.0234375,0.03125,0.0,-0.03125,-0.0078125,-0.015625,-0.046875,0.046875,-0.0,-0.0390625,-0.0546875,0.0078125,-0.03125,-0.015625,-0.0078125,-0.0078125,-0.0,-0.0078125,-0.015625,0.0234375,0.0234375,-0.0546875,-0.0234375,-0.015625,0.015625,-0.0,-0.0,-0.0234375,-0.03125,0.015625,-0.0078125,0.0703125,0.1328125,-0.0546875,0.015625,-0.03125,-0.0078125,0.0703125,0.0234375,-0.0078125,0.0078125,0.0078125,0.0,-0.0078125,-0.0,-0.015625,0.0,-0.0078125,-0.0078125,-0.0703125,-0.046875,-0.0390625,0.046875,0.0,0.03125,0.0546875,-0.0234375,-0.0234375,-0.015625,0.015625,-0.0078125,-0.015625,-0.0234375,-0.015625,0.0703125,0.046875,0.0078125,-0.0390625,-0.0546875,-0.0234375,0.0234375,-0.046875,0.0,0.0078125,0.03125,0.015625,0.0078125,0.015625,0.0,-0.0078125,-0.0,-0.0078125,0.0078125,0.0,-0.0234375,-0.0546875,-0.0078125,-0.0,-0.0390625,-0.046875,-0.0234375,0.015625,0.03125,-0.0,-0.0390625,0.125,-0.015625,-0.1015625,-0.015625,0.0,-0.015625,0.0234375,-0.0078125,-0.0234375,-0.046875,-0.0234375,0.03125,0.0390625,-0.0546875,0.0078125,-0.046875,-0.0078125,-0.0390625,0.015625,-0.0625,0.0625,0.0390625,0.015625,-0.015625,-0.015625,-0.015625,-0.03125,0.0,0.0390625,-0.015625,-0.03125,-0.0390625,0.0625,-0.0078125,-0.0078125,0.015625,-0.015625,-0.0,-0.03125,-0.0234375,-0.0234375,-0.0546875,-0.0234375,-0.0078125,-0.03125,-0.0,-0.0,0.015625,0.0,0.0078125,-0.0,0.0,0.0078125,0.0078125,0.0078125,0.0078125,-0.0078125,-0.0234375,0.0,0.0390625,0.09375,-0.0234375,-0.0078125,0.0390625,-0.0390625,0.015625,-0.0625,-0.015625,-0.0546875,0.140625,0.0,-0.078125,-0.0546875,-0.0703125,-0.0625,0.0234375,0.0234375,0.0625,-0.0078125,-0.0,-0.015625,-0.015625,0.0,-0.0078125,-0.015625,0.0078125,-0.0078125,0.015625,-0.0,0.0078125,0.0234375,0.0078125,-0.015625,-0.03125,-0.0390625,0.0078125,-0.0234375,-0.015625,-0.046875,-0.0859375,-0.046875,0.0390625,-0.03125,-0.0234375,-0.015625,-0.015625,-0.015625,0.015625,-0.0234375,-0.0078125,-0.015625,-0.0703125,0.015625,-0.0703125,0.0859375,0.015625,0.03125,-0.1171875,-0.0546875,0.0,-0.046875,-0.0078125,0.0234375,0.1796875,-0.0078125,-0.0,0.0390625,-0.0546875,0.0390625,-0.0546875,-0.03125,0.0078125,-0.046875,-0.0078125,0.03125,-0.0625,-0.0234375,0.0,-0.0859375,-0.0078125,-0.0078125,-0.0234375,-0.0078125,-0.0625,0.015625,-0.015625,-0.03125,0.046875,0.0078125,-0.0390625,-0.1484375,-0.0078125,0.0234375,-0.0078125,-0.0546875,0.0078125,-0.0625,-0.0625,-0.03125,0.0078125,-0.0078125,0.03125,-0.0390625,0.0,-0.0625,-0.0703125,-0.0078125,-0.03125,-0.0,0.015625,-0.046875,0.03125,0.015625,-0.015625,-0.0234375,-0.0,0.0234375,0.0234375,-0.0234375,-0.1171875,-0.0625,-0.0234375,0.1328125,0.046875,0.015625,0.0625,0.0078125,-0.015625,-0.0625,-0.0390625,-0.0,-0.046875,0.015625,0.015625,-0.0546875,-0.0234375,-0.0078125,-0.0234375,-0.078125,0.0390625,-0.03125,-0.0078125,0.0234375,-0.0390625,-0.109375,-0.0078125,-0.015625,-0.046875,0.046875,-0.0078125,-0.03125,0.0078125,0.015625,0.0625,-0.0234375,0.03125,0.09375,-0.0078125,0.0,0.0703125,0.0078125,-0.015625,-0.0859375,0.03125,0.0078125,-0.0390625,-0.0078125,-0.0234375,-0.0234375,0.03125,-0.046875,-0.0234375,-0.015625,-0.0078125,0.0234375,0.0,0.015625,0.015625,-0.0078125,-0.0078125,-0.0078125,-0.1015625,-0.015625,-0.0625,0.015625,-0.0390625,-0.0390625,0.03125,0.015625,-0.0,-0.0625,-0.0078125,-0.03125,-0.0078125,0.0859375,-0.0703125,0.03125,0.0078125,0.0234375,-0.0234375,-0.0703125,-0.046875,0.078125,-0.015625,0.0,-0.0625,-0.0546875,0.0,0.015625,0.0078125,-0.0078125,0.015625,0.0078125,-0.0078125,-0.0078125,0.0078125,0.0078125,-0.09375,0.1171875,-0.015625,0.0078125,-0.078125,-0.0390625,0.046875,-0.0078125,-0.015625,-0.0078125,-0.0078125,-0.0234375,-0.0078125,0.03125,-0.0078125,-0.046875,-0.0234375,-0.0,0.0625,-0.0390625,-0.0078125,-0.078125,-0.0,-0.03125,-0.0078125,-0.015625,-0.015625,-0.015625,-0.046875,-0.0078125,0.0078125,0.0625,0.0234375,0.015625,-0.03125,-0.015625,-0.046875,-0.0546875,0.03125,0.046875,-0.03125,0.015625,0.078125,0.046875,-0.03125,-0.0078125,0.0703125,0.0078125,0.015625,0.03125,0.0234375,-0.0078125,0.03125,-0.015625,0.0390625,-0.0234375,-0.0078125,0.015625,0.0,-0.0078125,0.0078125,0.0078125,0.0078125,0.015625,0.0,-0.015625,0.03125,0.0,-0.03125,0.0,-0.015625,-0.0,-0.015625,0.046875,0.015625,0.046875,-0.0,0.0234375,0.046875,-0.0546875,-0.046875,0.03125,-0.03125,-0.0390625,0.0078125,-0.0703125,0.03125,-0.046875,-0.0625,-0.0234375,0.0078125,0.0078125,0.0,0.0078125,0.0078125,0.0078125,0.0078125,-0.015625,0.0,0.03125,0.1015625,0.0390625,-0.03125,-0.0234375,0.0234375,-0.0078125,0.0,-0.0,0.0,-0.0078125,0.0546875,-0.015625,0.0390625,0.015625,-0.0234375,-0.0078125,-0.0234375,-0.03125,0.0,0.0390625,-0.0078125,-0.0625,0.1015625,-0.0,-0.0234375,-0.03125,0.0,0.046875,-0.0,-0.0625,-0.03125,0.03125,-0.0078125,-0.0546875,-0.0234375,0.046875,-0.0703125,-0.015625,0.03125,0.0234375,0.0703125,-0.015625,-0.03125,0.03125,-0.03125,0.015625,0.046875,0.0078125,-0.0546875,-0.0078125,0.0078125,-0.0625,-0.0,0.109375,-0.0390625,-0.0,-0.0703125,-0.0078125,0.0078125,0.03125,-0.015625,-0.0078125,0.0390625,-0.0,0.0390625,0.0703125,-0.046875,0.0078125,0.0,-0.0234375,-0.015625,0.0,0.0078125,0.03125,-0.015625,-0.0078125,-0.0390625,-0.0078125,-0.0390625,0.046875,0.0,-0.0703125,-0.03125,-0.0234375,-0.015625,-0.0234375,-0.046875,-0.0,-0.03125,0.046875,0.015625,-0.09375,0.03125,-0.015625,-0.046875,0.0078125,0.046875,-0.03125,-0.078125,-0.0234375,0.0390625,0.0234375,-0.0234375,-0.03125,0.0390625,-0.0,-0.015625,0.0234375,-0.0546875,0.0,0.0078125,-0.078125,-0.0234375,0.0859375,0.015625,0.0625,0.0,0.0,0.078125,-0.015625,-0.0546875,0.0,-0.015625,-0.0390625,-0.0234375,0.046875,0.0078125,-0.015625,-0.078125,-0.0390625,0.078125,-0.0234375,-0.046875,-0.015625,-0.0234375,0.0390625,0.0078125,0.0703125,0.0859375,0.0390625,-0.015625,-0.0546875,-0.0234375,0.0,-0.0078125,-0.0078125,0.0234375,-0.0078125,-0.0,-0.015625,-0.0078125,0.0078125,-0.0078125,0.078125,-0.015625,0.078125,0.015625,0.046875,0.03125,-0.03125,-0.0625,-0.015625,-0.015625,-0.0234375,-0.0078125,-0.0078125,-0.078125,0.0078125,0.0390625,0.1953125,-0.0078125,-0.0703125,-0.046875,-0.015625,-0.046875,-0.046875,-0.0234375,0.078125,0.140625,-0.0078125,0.0078125,-0.0078125,0.0078125,0.0,0.0,0.0,-0.0,-0.0,-0.03125,-0.0859375,-0.1015625,-0.046875,-0.0625,0.0234375,0.03125,0.09375,0.0625,-0.0390625,-0.0625,0.046875,-0.0,0.0546875,0.0234375,-0.015625,-0.0859375,-0.0078125,-0.03125,-0.0234375,-0.0234375,-0.1015625,0.0078125,-0.1484375,-0.0390625,-0.0078125,0.0234375,-0.0390625,-0.046875,-0.046875,-0.0078125,-0.0625,-0.0390625,0.0703125,-0.015625,0.0234375,-0.015625,-0.0625,-0.0234375,0.015625,0.0546875,-0.0078125,-0.0703125,0.0546875,0.03125,-0.015625,-0.0078125,0.0234375,0.0078125,-0.0234375,0.0625,0.0625,0.0703125,0.0390625,0.015625,0.015625,-0.015625,0.015625,0.0546875,0.0390625,-0.0390625,0.0078125,-0.0625,-0.015625,-0.03125,-0.0234375,-0.0390625,-0.0,-0.0390625,0.0390625,0.0,-0.0078125,-0.03125,-0.015625,-0.0546875,0.0390625,-0.1171875,-0.078125,-0.0078125,0.15625,-0.046875,-0.0390625,-0.0234375,-0.03125,0.0625,-0.0859375,0.0703125,0.0234375,-0.0703125,-0.015625,-0.0078125,-0.0078125,0.0078125,-0.0,-0.0078125,-0.015625,0.0078125,0.0,-0.0,-0.0390625,-0.046875,-0.0078125,0.0234375,0.046875,-0.03125,-0.0,-0.0390625,-0.0703125,0.046875,0.015625,0.015625,0.0,-0.046875,0.0234375,-0.0078125,-0.078125,0.09375,-0.0390625,-0.046875,-0.0234375,0.0546875,-0.0,-0.0234375,0.03125,0.0234375,-0.015625,-0.03125,0.0,-0.0234375,0.0390625,-0.046875,0.109375,0.0234375,-0.0390625,0.0078125,0.0234375,-0.0390625,-0.0234375,-0.0625,-0.015625,-0.0,0.03125,-0.03125,0.0390625,0.03125,0.0390625,0.0234375,0.078125,-0.09375,0.03125,0.0234375,-0.046875,0.0234375,-0.0078125,-0.0859375,-0.0234375,-0.1015625,0.0390625,-0.109375,0.0390625,0.0234375,0.0625,-0.046875,-0.03125,-0.015625,0.0703125,0.0859375,-0.0625,0.03125,0.0859375,0.0625,0.0,0.0625,0.0390625,-0.0390625,-0.015625,0.0078125,-0.09375,0.0078125,-0.140625,0.046875,-0.0078125,0.0,-0.0390625,0.03125,-0.03125,-0.03125,0.0078125,-0.0078125,-0.015625,-0.03125,-0.015625,-0.1484375,-0.0546875,-0.015625,-0.0234375,0.1015625,-0.1171875,0.0078125,-0.0078125,-0.03125,-0.046875,-0.1875,-0.015625,-0.0625,0.109375,-0.0546875,0.03125,-0.0390625,0.046875,-0.0234375,0.0078125,0.0078125,-0.078125,0.015625,-0.109375,-0.03125,0.0390625,-0.03125,0.0546875,-0.1015625,0.015625,0.0703125,0.0,-0.03125,0.015625,-0.0390625,0.046875,-0.0390625,0.0546875,-0.0625,0.0546875,0.0,-0.0390625,0.0390625,0.0703125,-0.015625,-0.0390625,-0.0703125,-0.0,-0.015625,-0.015625,0.0,-0.0078125,-0.0,-0.015625,-0.0078125,0.015625,-0.0078125,-0.0,0.015625,0.0078125,-0.0234375,-0.109375,-0.1015625,-0.0078125,0.0234375,-0.0078125,0.0234375,-0.015625,0.0234375,0.046875,0.015625,0.0390625,-0.0390625,0.1015625,0.0078125,0.0234375,-0.046875,0.0625,-0.0078125,0.0390625,0.125,0.0,-0.109375,0.0078125,0.0390625,-0.03125,-0.0078125,-0.0078125,0.0078125,-0.0,-0.0078125,0.0078125,0.0,0.0078125,0.0078125,-0.015625,-0.0703125,-0.015625,0.078125,-0.0546875,-0.0078125,0.0390625,-0.0,-0.0625,-0.015625,-0.0078125,-0.0859375,-0.0234375,0.15625,0.0078125,0.078125,0.0390625,0.03125,0.03125,0.0234375,-0.1171875,0.0078125,-0.0078125,0.0078125,0.0390625,-0.0078125,-0.0078125,0.0078125,-0.0703125,-0.0703125,-0.0234375,0.03125,0.0234375,0.0,-0.0078125,0.03125,0.015625,-0.0625,0.0546875,-0.0,0.0,-0.0390625,0.0234375,-0.0390625,0.015625,-0.0078125,-0.0078125,0.0078125,-0.0078125,-0.0390625,-0.015625,-0.0234375,0.015625,0.0078125,0.0234375,-0.015625,-0.015625,-0.0078125,0.0078125,0.03125,-0.015625,0.0078125,0.0078125,0.0234375,0.0234375,-0.0546875,0.046875,0.03125,0.03125,-0.09375,0.0078125,0.0078125,0.015625,0.0859375,-0.0078125,0.015625,-0.015625,0.0,0.03125,-0.09375,0.0078125,0.015625,-0.0234375,0.015625,-0.046875,0.0234375,0.078125,-0.0234375,0.0,-0.0078125,-0.015625,0.0,-0.0234375,0.0234375,0.0,0.0234375,-0.0,0.0078125,0.0,-0.0078125,-0.0078125,0.015625,-0.046875,-0.0078125,0.0078125,-0.0234375,-0.015625,-0.0234375,-0.015625,0.0234375,0.0,0.0546875,0.0078125,-0.0390625,-0.0546875,0.0234375,0.0078125,0.015625,-0.0078125,-0.0625,-0.03125,0.015625,0.046875,0.046875,-0.0078125,-0.0390625,0.015625,-0.046875,-0.0234375,0.0234375,0.0078125,-0.015625,-0.0625,0.03125,-0.0390625,-0.015625,0.0234375,0.0234375,0.015625,0.015625,0.046875,-0.0390625,-0.0625,-0.0703125,-0.0078125,0.0078125,-0.0703125,0.0,0.0078125,-0.0546875,0.0234375,0.015625,-0.03125,-0.046875,0.0703125,-0.0078125,0.0703125,-0.0546875,-0.046875,-0.0546875,-0.03125,-0.0390625,0.0078125,-0.0390625,0.015625,-0.0,-0.0234375,-0.015625,-0.015625,-0.0078125,-0.046875,-0.0390625,0.0390625,0.0390625,0.046875,-0.046875,-0.0234375,0.0546875,0.0078125,0.0234375,-0.0,0.0078125,-0.03125,-0.015625,-0.0078125,0.078125,0.046875,0.0234375,-0.046875,0.0703125,0.0,-0.0234375,0.015625,-0.1171875,0.03125,-0.0625,-0.0234375,-0.0390625,-0.0546875,-0.0,0.125,0.03125,0.078125,-0.0859375,0.0078125,0.0,-0.0,0.0078125,0.046875,-0.1171875,0.03125,0.0390625,-0.015625,0.109375,-0.0234375,-0.0234375,-0.0078125,-0.078125,0.0234375,0.03125,-0.0,-0.0234375,-0.015625,0.0390625,0.03125,-0.0078125,0.1171875,-0.078125,-0.015625,0.0703125,-0.0546875,-0.0703125,-0.015625,-0.015625,0.0234375,-0.0234375,0.0078125,-0.0390625,0.0625,-0.0546875,0.0625,-0.0703125,0.0078125,-0.03125,0.0,0.0,-0.0,0.0078125,-0.015625,-0.015625,-0.0078125,-0.015625,-0.0234375,0.0078125,0.0625,0.0625,-0.0234375,0.0,-0.0546875,-0.0234375,-0.0,-0.0078125,-0.0078125,-0.0078125,-0.0078125,-0.0078125,-0.046875,-0.0859375,0.046875,0.0078125,0.09375,0.0078125,-0.0625,0.109375,0.046875,0.0,-0.0546875,0.0,-0.0546875,0.078125,0.0078125,0.0234375,0.0078125,-0.0078125,0.0,0.0078125,0.0,-0.0078125,-0.015625,0.0703125,0.0703125,0.0390625,0.046875,-0.0859375,-0.0234375,0.09375,-0.0234375,0.03125,-0.0078125,-0.0,-0.03125,-0.125,-0.078125,-0.078125,0.0234375,-0.0,-0.0234375,0.0546875,-0.078125,0.015625,0.015625,-0.0703125,0.0078125,0.078125,-0.046875,0.0234375,-0.015625,0.0546875,-0.03125,-0.0,-0.03125,0.03125,0.0078125,0.0625,0.015625,-0.0390625,0.0234375,-0.015625,0.0546875,-0.0234375,-0.0390625,0.0625,0.0,0.125,-0.0078125,-0.0078125,-0.0390625,0.046875,-0.0078125,-0.0078125,0.015625,-0.0390625,-0.046875,-0.0078125,-0.078125,-0.015625,0.0078125,0.046875,0.015625,0.0078125,0.015625,-0.0078125,0.0,0.0390625,-0.0234375,0.03125,-0.015625,-0.0078125,0.015625,0.0546875,-0.03125,0.0078125,-0.015625,0.0390625,0.046875,0.0390625,0.046875,-0.0078125,-0.0546875,-0.0078125,0.0,-0.03125,-0.0234375,-0.046875,0.1015625,-0.0234375,0.015625,0.0546875,-0.015625,-0.015625,-0.015625,-0.0078125,-0.03125,-0.0078125,-0.015625,0.0,0.0234375,-0.0078125,-0.015625,0.03125,0.015625,-0.0390625,0.0078125,-0.0078125,0.0,-0.0,-0.0078125,-0.078125,-0.0,0.0078125,-0.078125,-0.0,0.046875,0.0234375,-0.0703125,-0.0078125,0.0234375,-0.0390625,-0.0078125,0.015625,0.0546875,0.046875,0.0234375,-0.09375,-0.046875,-0.0625,0.0234375,-0.03125,-0.046875,-0.03125,-0.0859375,-0.0078125,0.0,-0.0,0.015625,-0.078125,-0.0078125,-0.0078125,-0.015625,0.0234375,0.0234375,0.046875,0.0859375,-0.0078125,0.0078125,-0.015625,0.0078125,-0.09375,0.03125,0.1015625,-0.046875,0.0234375,-0.078125,-0.09375,-0.046875,-0.0859375,0.0390625,-0.09375,0.15625,-0.0390625,0.0703125,-0.078125,0.0078125,-0.015625,0.046875,-0.0546875,-0.03125,0.0390625,-0.046875,0.0390625,-0.078125,-0.03125,-0.0234375,-0.03125,-0.0859375,-0.015625,0.0546875,0.0546875,0.0390625,-0.0,0.03125,0.0390625,0.0,-0.0234375,-0.0390625,0.0078125,-0.015625,-0.0,0.0859375,-0.0078125,-0.078125,-0.0703125,0.015625,-0.0703125,-0.015625,0.1484375,-0.0078125,-0.0390625,-0.03125,0.0,0.0390625,0.0546875,-0.0,-0.0,0.0,0.0078125,0.0234375,-0.0390625,-0.0078125,0.0,-0.1015625,-0.0625,0.234375,-0.046875,0.2109375,0.0078125,0.1171875,-0.0390625,-0.046875,-0.0234375,-0.015625,0.0078125,-0.1171875,0.0234375,-0.0546875,-0.046875,-0.109375,0.0703125,-0.0546875,0.03125,0.03125,0.0078125,-0.0546875,-0.0234375,-0.0390625,-0.046875,-0.015625,0.03125,0.03125,-0.015625,-0.0546875,-0.0390625,-0.0234375,-0.0078125,-0.0078125,0.0,0.0078125,-0.015625,0.0078125,0.015625,0.0078125,0.0234375,-0.046875,-0.0234375,-0.0,0.0,0.015625,-0.015625,-0.0234375,-0.046875,0.0703125,0.03125,0.0234375,-0.015625,-0.0234375,-0.015625,-0.0078125,-0.03125,-0.0078125,-0.078125,0.109375,-0.0234375,-0.0234375,-0.0078125,-0.0234375,0.015625,0.0234375,-0.0078125,0.0078125,-0.0078125,0.015625,-0.0078125,-0.0078125,-0.0078125,0.0078125,-0.0078125,0.0,0.0703125,-0.046875,0.0,0.015625,-0.046875,-0.015625,0.015625,-0.0,-0.046875,0.0390625,0.0078125,-0.015625,0.046875,-0.0234375,0.046875,-0.0078125,0.015625,0.0234375,0.09375,-0.0859375,-0.0390625,0.015625,-0.0234375,0.0078125,0.015625,-0.0390625,-0.0078125,0.046875,-0.0078125,-0.0078125,-0.0234375,-0.0546875,0.0,0.0,-0.03125,-0.0,-0.015625,-0.015625,0.015625,-0.0078125,-0.0390625,-0.0625,0.046875,0.015625,0.03125,-0.0546875,0.0234375,0.015625,0.0078125,0.0078125,0.015625,0.015625,0.0078125,-0.0,0.0078125,-0.015625,-0.03125,-0.0078125,0.0234375,-0.0,0.0078125,0.0078125,0.0078125,-0.0078125,0.03125,-0.0078125,0.046875,-0.0078125,-0.0234375,-0.015625,0.0,0.015625,-0.015625,-0.0859375,0.0078125,-0.0390625,-0.0234375,-0.0,-0.0234375,-0.0390625,-0.0234375,-0.0078125,-0.078125,-0.0625,0.0625,0.0078125,-0.015625,-0.0078125,-0.0078125,-0.0,-0.0078125,-0.0078125,0.0078125,-0.015625,-0.0078125,-0.0078125,-0.0078125,0.0,0.0,-0.0,-0.015625,-0.0234375,-0.015625,-0.0078125,0.0,0.015625,-0.0234375,0.0078125,0.0234375,0.0625,0.046875,-0.0078125,0.0078125,-0.0234375,0.0078125,-0.0546875,0.0,-0.0859375,-0.015625,-0.015625,-0.0,0.0234375,0.0,-0.0234375,0.0078125,-0.0234375,-0.03125,-0.0078125,0.078125,0.015625,0.046875,-0.03125,0.0078125,0.03125,0.0234375,-0.0390625,0.0625,-0.03125,-0.015625,-0.0234375,-0.046875,-0.0234375,-0.0390625,-0.0234375,-0.078125,-0.0078125,0.0078125,0.03125,0.0078125,-0.0859375,-0.015625,-0.0234375,-0.0234375,-0.0546875,0.0859375,0.109375,0.03125,-0.03125,-0.0234375,-0.0546875,-0.0078125,0.0078125,-0.046875,-0.0,-0.015625,-0.03125,0.0234375,-0.078125,0.0078125,0.0234375,-0.0234375,0.0078125,-0.015625,0.0234375,0.0234375,-0.0234375,0.046875,0.0234375,-0.0234375,0.015625,0.0234375,0.0390625,0.0078125,-0.0625,-0.0078125,0.0,-0.015625,0.03125,0.0078125,0.0234375,-0.046875,0.0625,0.015625,-0.0390625,0.0078125,-0.0078125,-0.0390625,0.03125,-0.03125,0.0078125,0.078125,-0.0234375,0.0,-0.09375,0.0078125,0.015625,0.015625,0.0703125,0.0234375,0.0,-0.015625,-0.046875,0.0078125,-0.046875,-0.0390625,-0.015625,-0.0078125,-0.015625,-0.0078125,0.03125,0.0390625,-0.0390625,-0.03125,0.0,-0.0078125,0.0078125,0.0859375,-0.0234375,0.0625,-0.0234375,-0.0390625,0.015625,-0.03125,-0.0,-0.0234375,0.0234375,-0.0390625,-0.0390625,-0.015625,-0.0546875,0.0625,0.015625,-0.03125,-0.015625,-0.015625,-0.015625,-0.0078125,0.0,-0.015625,0.0,0.0078125,0.0078125,-0.0,-0.09375,-0.0078125,-0.0390625,-0.09375,-0.015625,-0.015625,0.0546875,0.0,0.0390625,-0.0390625,-0.0078125,0.078125,-0.015625,0.0234375,0.0546875,-0.0390625,-0.0078125,-0.078125,-0.046875,-0.0625,0.0078125,-0.078125,-0.0234375,0.015625,-0.0703125,0.015625,-0.0,-0.015625,-0.0,-0.015625,0.015625,-0.0,0.0,0.0,-0.0078125,-0.0078125,-0.09375,-0.0234375,0.046875,-0.0,0.109375,0.015625,0.0,0.015625,-0.0078125,0.046875,-0.03125,-0.1015625,0.0078125,-0.0390625,0.03125,0.0625,0.0,-0.03125,-0.0546875,-0.0234375,-0.0703125,-0.0,-0.015625,0.1171875,0.0859375,-0.046875,-0.0078125,-0.0703125,0.0078125,-0.0390625,0.03125,0.0,-0.03125,0.0390625,-0.0390625,-0.0078125,0.046875,-0.03125,0.046875,0.0078125,0.03125,0.0703125,-0.0390625,0.0234375,-0.015625,0.015625,0.0,-0.0546875,-0.0546875,-0.0390625,-0.0390625,-0.0078125,0.0234375,0.0234375,-0.03125,0.0078125,-0.0390625,0.0234375,-0.0390625,-0.0234375,-0.0078125,0.0078125,-0.015625,-0.0078125,-0.0234375,0.0390625,-0.0078125,-0.0,0.0078125,0.0390625,-0.03125,-0.0234375,0.0703125,0.0390625,-0.0625,0.0546875,-0.0625,0.1171875,0.0078125,-0.0234375,0.0078125,-0.078125,0.046875,0.046875,-0.03125,0.0234375,0.0234375,0.0390625,0.0859375,0.015625,-0.0078125,-0.0078125,0.015625,0.0234375,0.0,0.0078125,0.0,-0.0078125,0.0546875,-0.0234375,0.0234375,-0.078125,-0.03125,-0.0078125,-0.0078125,-0.0234375,0.0078125,0.03125,0.0625,0.0,0.0625,0.0078125,-0.0546875,-0.015625,-0.0078125,-0.0234375,-0.046875,0.015625,-0.015625,-0.0078125,0.03125,-0.0703125,-0.046875,0.046875,-0.0390625,0.0078125,0.0234375,-0.03125,-0.03125,0.1640625,-0.0234375,-0.015625,0.0078125,-0.0390625,0.0,-0.03125,0.0390625,-0.015625,0.03125,0.0078125,0.03125,-0.078125,0.03125,0.0703125,-0.0078125,0.109375,0.0234375,-0.03125,0.0,-0.015625,-0.0,-0.0078125,0.0234375,-0.015625,-0.0234375,-0.0859375,-0.0859375,-0.0703125,-0.015625,0.0390625,-0.0078125,0.0078125,-0.0390625,0.0078125,-0.0390625,-0.046875,-0.0703125,0.0078125,-0.0859375,-0.0078125,0.0390625,0.0234375,0.0234375,-0.0703125,0.0390625,-0.1015625,-0.0546875,0.0,-0.1015625,0.0234375,-0.0546875,-0.0078125,-0.03125,0.0390625,-0.0390625,-0.0078125,0.0078125,0.0234375,0.1328125,-0.140625,0.015625,0.0546875,-0.03125,0.0234375,-0.0234375,-0.125,-0.0234375,-0.0390625,-0.109375,-0.0859375,0.078125,-0.015625,-0.046875,0.078125,0.203125,0.03125,0.0234375,-0.1015625,-0.0625,-0.0,0.03125,-0.015625,-0.0546875,0.0546875,0.0078125,0.0078125,0.03125,0.015625,-0.0546875,-0.0,-0.03125,-0.0625,0.0703125,-0.0078125,0.1015625,-0.015625,0.0,0.0390625,0.0,0.03125,-0.0,-0.0546875,0.0,0.0390625,0.03125,-0.0078125,-0.0078125,0.015625,-0.0078125,-0.0,0.0234375,-0.0,-0.0078125,-0.0078125,0.015625,0.0078125,0.015625,-0.0078125,-0.0078125,0.0,-0.0078125,0.1640625,-0.0,0.015625,0.078125,-0.0546875,0.0078125,-0.0078125,0.0078125,0.03125,-0.0,0.015625,0.0390625,0.015625,-0.0234375,-0.015625,-0.0078125,-0.0390625,-0.0,0.0078125,-0.03125,0.0234375,0.0625,-0.015625,-0.0234375,-0.0625,-0.0234375,0.0078125,-0.015625,-0.0078125,0.0078125,-0.0078125,0.0078125,-0.015625,-0.015625,0.015625,-0.0,0.0390625,0.0546875,0.0078125,0.0390625,-0.0390625,-0.0703125,-0.015625,0.0,-0.0078125,-0.0078125,0.015625,-0.0234375,-0.03125,0.0234375,-0.0390625,-0.03125,-0.03125,0.03125,0.0078125,-0.09375,0.015625,0.0546875,-0.015625,0.0078125,0.0,-0.015625,-0.0078125,0.015625,-0.015625,0.0078125,-0.03125,0.0078125,0.0,0.0078125,-0.0078125,-0.0078125,0.0,0.0625,-0.046875,-0.015625,0.09375,-0.0234375,-0.0390625,-0.0234375,-0.0,-0.0078125,0.03125,-0.0078125,-0.0078125,0.0078125,-0.015625,0.015625,0.0390625,0.0,-0.03125,0.0,-0.0078125,-0.0390625,-0.0078125,-0.015625,-0.0078125,-0.0,0.0234375,-0.015625,0.0078125,0.0078125,-0.03125,-0.046875,0.046875,0.0234375,-0.0,-0.0,-0.015625,-0.0,-0.0390625,-0.0703125,0.0078125,-0.0078125,-0.0,-0.0234375,0.0078125,0.078125,0.0234375,-0.0078125,-0.046875,0.0234375,0.0078125,-0.0078125,-0.046875,0.015625,0.015625,0.0390625,0.0,0.0,-0.0234375,-0.0078125,-0.015625,0.0078125,-0.015625,0.03125,-0.03125,-0.0078125,0.015625,0.015625,-0.03125,-0.0078125,0.015625,-0.015625,-0.015625,-0.046875,0.0078125,-0.0234375,0.015625,0.0078125,0.0234375,-0.0234375,-0.0078125,0.0703125,0.0,0.03125,-0.0859375,0.015625,-0.0546875,-0.0,-0.0,0.015625,0.0390625,0.09375,0.03125,-0.015625,-0.0625,-0.0078125,-0.0703125,-0.0546875,0.0234375,0.0703125,0.0859375,-0.046875,-0.0625,-0.03125,-0.0234375,-0.0625,-0.0546875,-0.03125,0.0234375,0.015625,-0.03125,0.015625,-0.0390625,0.0078125,-0.015625,-0.0078125,0.0,0.015625,-0.0625,-0.0078125,0.09375,-0.0625,0.0390625,-0.03125,-0.0390625,0.0234375,-0.0078125,-0.046875,-0.015625,-0.0,-0.0234375,0.0078125,0.015625,0.015625,-0.0234375,-0.0859375,-0.015625,0.046875,-0.0390625,-0.0,0.015625,-0.0,0.0234375,0.015625,0.0703125,0.078125,0.0390625,0.0078125,-0.046875,-0.0078125,-0.0234375,-0.0234375,0.0,-0.1015625,-0.0234375,-0.015625,-0.0625,-0.0234375,0.0390625,-0.0078125,0.046875,0.015625,0.03125,0.03125,0.0078125,0.0,-0.0546875,0.0078125,-0.0390625,-0.03125,0.015625,0.046875,0.0234375,0.015625,0.03125,-0.0078125,0.0078125,0.0390625,-0.0625,-0.0234375,0.0859375,0.0,0.015625,0.0078125,-0.03125,-0.015625,-0.015625,-0.015625,0.0,-0.0234375,0.03125,-0.0390625,-0.078125,0.0234375,-0.0,-0.03125,-0.03125,0.0,0.046875,0.0546875,-0.03125,-0.078125,0.09375,-0.0859375,0.0078125,-0.0234375,0.046875,0.0078125,0.0,0.015625,0.0078125,-0.0,-0.0234375,-0.015625,0.0078125,0.0,-0.0234375,-0.0,0.0,-0.0078125,0.015625,0.0234375,0.0,-0.03125,0.015625,-0.03125,-0.0078125,0.0546875,0.03125,-0.015625,-0.03125,0.0234375,-0.0234375,-0.015625,-0.0625,-0.0078125,-0.046875,0.015625,0.0234375,-0.015625,-0.015625,-0.03125,-0.0078125,-0.0,-0.015625,-0.0,0.0078125,0.0078125,-0.0078125,0.0078125,-0.0078125,0.0,-0.0234375,-0.015625,-0.015625,0.0703125,-0.09375,-0.1015625,0.015625,-0.0234375,-0.0546875,0.0546875,0.0078125,0.0390625,-0.0546875,0.0078125,-0.015625,0.046875,-0.0078125,0.0234375,0.0234375,0.0234375,-0.03125,-0.0390625,-0.078125,-0.046875,-0.0859375,-0.0,0.046875,0.015625,-0.125,-0.046875,-0.0546875,0.03125,0.1015625,-0.046875,-0.0234375,0.0546875,-0.0234375,-0.0078125,-0.0234375,0.0390625,0.0078125,0.0546875,0.0703125,-0.0,0.0625,0.0390625,0.0234375,-0.015625,-0.03125,-0.0234375,-0.03125,-0.046875,-0.015625,-0.0078125,0.0234375,0.0390625,0.046875,-0.0078125,-0.0078125,0.015625,-0.015625,-0.0,-0.015625,-0.015625,0.0390625,0.03125,-0.0234375,-0.015625,-0.0234375,0.0,0.09375,-0.0390625,0.078125,-0.03125,0.0390625,-0.0234375,-0.046875,-0.0234375,0.015625,0.0234375,0.1015625,0.0078125,-0.046875,-0.1015625,0.0625,-0.0390625,0.015625,-0.03125,-0.0234375,0.0390625,-0.0,-0.015625,-0.0078125,0.0234375,0.0234375,0.0234375,0.0234375,0.0078125,0.0234375,0.015625,-0.0234375,-0.0078125,-0.0234375,-0.015625,-0.015625,0.0078125,-0.0078125,-0.0234375,0.0234375,-0.0,0.1171875,0.0390625,-0.0546875,-0.046875,0.0390625,0.0390625,0.03125,0.0,0.0078125,0.0234375,-0.078125,0.0,0.015625,-0.0703125,-0.0625,-0.046875,0.046875,-0.09375,0.046875,-0.0078125,0.0234375,0.0390625,-0.0546875,0.0234375,0.015625,0.0390625,0.03125,0.0078125,-0.0234375,-0.0390625,-0.015625,0.0546875,-0.125,0.0,0.0390625,0.0234375,0.0703125,-0.0234375,-0.0078125,-0.046875,-0.0078125,0.0234375,0.0234375,0.0625,0.0546875,0.046875,-0.03125,-0.0703125,-0.0078125,-0.0390625,0.015625,-0.0234375,-0.0078125,0.0234375,0.015625,-0.0625,0.03125,-0.0078125,0.0078125,-0.0625,0.046875,0.0390625,0.0234375,0.0703125,-0.0078125,0.046875,-0.0703125,0.0234375,-0.015625,0.09375,0.046875,0.046875,0.0859375,-0.0078125,-0.0234375,-0.015625,0.0234375,0.0625,-0.078125,-0.03125,-0.0703125,0.015625,0.0546875,-0.078125,0.0625,0.0078125,0.03125,0.03125,-0.0078125,-0.0546875,-0.046875,-0.0078125,-0.0546875,0.03125,0.0234375,0.1015625,0.0703125,0.03125,-0.0,0.03125,-0.0234375,0.03125,0.0703125,-0.0078125,0.03125,0.015625,-0.03125,-0.0078125,0.046875,-0.0625,0.0390625,-0.0078125,0.0,0.0234375,-0.0234375,0.0625,0.0546875,0.0703125,0.0078125,-0.0546875,-0.0546875,-0.09375,-0.1171875,-0.046875,0.0,0.015625,0.0078125,0.0078125,-0.03125,0.015625,-0.015625,0.046875,0.0859375,0.015625,-0.0078125,0.0078125,-0.0078125,-0.0078125,0.0234375,-0.0,0.0078125,-0.0078125,0.0,-0.0078125,0.015625,0.0078125,0.015625,-0.03125,-0.0859375,0.0,-0.0234375,0.0078125,-0.0078125,0.015625,0.09375,-0.046875,0.0546875,0.0,-0.015625,0.0234375,-0.0078125,0.0234375,-0.0,-0.0078125,0.0390625,-0.015625,-0.015625,-0.0625,-0.03125,-0.0078125,-0.0078125,0.0078125,-0.015625,-0.015625,-0.015625,-0.0,0.0,0.0078125,-0.0234375,-0.0234375,-0.0234375,0.0078125,-0.09375,-0.046875,0.1015625,-0.0703125,0.0078125,-0.0078125,-0.0390625,-0.0078125,-0.1015625,0.0,-0.0,0.1171875,0.0703125,0.0703125,-0.015625,-0.0234375,0.0,0.0078125,-0.0234375,0.0078125,-0.015625,-0.0546875,-0.03125,0.0078125,-0.0078125,-0.03125,-0.0234375,0.0625,0.015625,0.0078125,0.0390625,0.03125,0.0078125,-0.046875,0.0078125,0.0234375,-0.015625,-0.0234375,-0.0390625,-0.015625,0.03125,-0.015625,-0.0234375,-0.0078125,0.015625,0.0078125,-0.0,-0.015625,-0.0234375,-0.0078125,-0.0078125,-0.0234375,-0.0078125,0.0078125,-0.0390625,0.015625,0.0234375,-0.015625,0.0078125,0.0390625,0.015625,-0.0078125,-0.0078125,0.046875,-0.0,-0.0234375,0.0234375,-0.0234375,0.03125,0.015625,0.0078125,-0.0703125,-0.0390625,-0.09375,0.171875,-0.1171875,0.0234375,-0.03125,-0.0078125,-0.015625,-0.0546875,-0.0546875,0.0,0.0546875,-0.109375,0.0625,0.015625,0.0234375,-0.0078125,-0.0078125,0.0078125,0.0,-0.0,0.0078125,0.0,0.0,-0.0078125,-0.0078125,0.015625,0.015625,-0.0078125,0.015625,0.0234375,-0.0234375,0.0234375,-0.0234375,-0.0234375,-0.03125,-0.0859375,0.015625,0.0390625,0.0390625,0.046875,-0.0234375,-0.0234375,-0.03125,-0.0703125,0.0078125,0.0078125,-0.03125,-0.0,0.0078125,0.03125,-0.0,-0.0546875,-0.140625,0.03125,-0.03125,-0.015625,0.0546875,0.0234375,-0.015625,-0.046875,-0.0390625,-0.0078125,-0.09375,-0.0078125,0.078125,-0.0234375,0.09375,-0.03125,-0.0234375,0.0078125,-0.015625,-0.0546875,0.078125,-0.0,-0.0390625,-0.0390625,-0.03125,-0.0078125,-0.015625,0.0546875,0.0078125,0.0390625,-0.0390625,-0.0625,-0.0234375,-0.0234375,-0.0,-0.015625,-0.0078125,0.0,-0.015625,-0.0546875,-0.046875,-0.0546875,0.0390625,0.0546875,0.015625,-0.015625,0.015625,-0.03125,0.03125,-0.0078125,0.0390625,-0.0078125,0.015625,0.0,0.0390625,0.0234375,0.09375,-0.0390625,0.0234375,0.0234375,-0.0,-0.03125,-0.0234375,0.0546875,-0.1015625,0.09375,0.046875,-0.046875,-0.0,0.0234375,0.0,-0.046875,-0.0703125,0.046875,-0.0078125,0.09375,0.03125,0.03125,0.0078125,-0.0234375,-0.0,0.078125,0.015625,0.0234375,-0.0625,-0.0390625,-0.015625,-0.0234375,-0.03125,-0.0078125,-0.0390625,0.1640625,-0.03125,0.03125,0.0078125,-0.03125,-0.0703125,-0.0234375,-0.0234375,0.1171875,-0.0625,0.046875,-0.0625,-0.0703125,-0.0078125,-0.046875,0.0,-0.0,-0.0390625,-0.015625,-0.0078125,-0.0234375,-0.0078125,0.0078125,0.015625,-0.0078125,-0.0078125,0.0234375,0.015625,-0.015625,-0.0078125,-0.0078125,0.0,-0.0078125,0.015625,0.0078125,0.0234375,-0.0234375,-0.0234375,0.03125,-0.015625,-0.0078125,-0.0234375,0.0546875,-0.0078125,-0.0078125,0.015625,-0.0,-0.015625,0.015625,0.0,-0.0546875,0.0390625,-0.0078125,-0.0,0.0078125,-0.015625,0.03125,0.0390625,-0.0234375,-0.0078125,-0.0,0.0078125,0.015625,-0.0078125,0.0078125,-0.0078125,-0.0078125,0.0,-0.0390625,0.0546875,-0.015625,-0.03125,0.0390625,-0.015625,0.078125,0.03125,-0.0,0.0390625,-0.046875,-0.0078125,0.03125,-0.0546875,-0.0234375,-0.046875,-0.0234375,-0.0078125,0.03125,0.0,-0.0078125,-0.09375,-0.0,-0.0,0.015625,-0.015625,-0.0078125,0.046875,-0.0234375,-0.0078125,0.0390625,0.0,-0.0234375,0.046875,0.015625,0.0,0.015625,-0.0390625,-0.015625,-0.0234375,-0.015625,-0.0,0.0234375,-0.03125,0.015625,-0.0625,-0.046875,0.0078125,-0.0,-0.0390625,0.0,0.0078125,-0.0078125,-0.015625,-0.015625,-0.0234375,-0.0,-0.0078125,0.0,-0.0078125,0.0,0.0078125,-0.015625,-0.03125,-0.0078125,0.0,-0.03125,0.015625,-0.015625,0.03125,-0.03125,-0.0,-0.0546875,-0.0546875,-0.0,0.078125,0.0078125,0.015625,-0.0625,-0.015625,-0.015625,0.046875,0.09375,-0.015625,-0.1015625,0.0390625,-0.015625,0.0078125,0.0390625,-0.015625,0.015625,0.0078125,-0.015625,-0.0078125,-0.0,-0.0,-0.0,-0.0078125,-0.0078125,-0.03125,-0.0546875,0.0078125,0.0078125,0.015625,-0.0078125,0.0078125,-0.0078125,0.0078125,-0.0,-0.0234375,0.0,0.0390625,-0.0859375,0.0,0.0625,0.0234375,-0.0078125,0.0703125,-0.046875,0.0,0.1484375,-0.078125,-0.0078125,-0.0234375,0.0078125,-0.0,-0.0546875,0.0078125,-0.015625,-0.015625,0.0078125,-0.03125,-0.046875,0.046875,-0.0,-0.0234375,-0.0234375,-0.0078125,-0.0546875,0.0390625,-0.0234375,0.0390625,0.0625,-0.0234375,-0.0546875,-0.0234375,-0.0078125,-0.0625,-0.03125,-0.0078125,-0.0390625,0.0234375,-0.0078125,-0.078125,-0.0078125,-0.0,0.078125,-0.0546875,-0.015625,-0.0234375,-0.0234375,0.0078125,0.03125,-0.0078125,-0.0,-0.0234375,0.046875,-0.0234375,-0.0390625,-0.015625,0.0,-0.03125,-0.0078125,0.0078125,-0.015625,-0.0234375,-0.0,-0.0234375,0.0078125,-0.015625,-0.015625,-0.0078125,-0.0078125,-0.03125,0.0078125,-0.015625,0.0390625,-0.0078125,-0.0078125,-0.015625,-0.0625,0.015625,-0.03125,0.015625,-0.0234375,0.0,-0.0546875,-0.0234375,0.015625,0.0859375,-0.0,0.09375,-0.0234375,-0.03125,-0.0625,-0.0078125,-0.0234375,-0.046875,0.0625,-0.0078125,0.015625,-0.015625,-0.0234375,0.015625,-0.078125,0.0,0.015625,-0.0,-0.0078125,0.046875,-0.0234375,-0.0078125,-0.015625,0.0234375,-0.0078125,-0.0625,-0.0546875,0.015625,0.0078125,-0.078125,-0.0234375,0.0,0.015625,-0.015625,-0.0234375,-0.015625,-0.0234375,0.03125,0.015625,0.046875,0.0078125,0.046875,-0.0390625,-0.0078125,-0.015625,0.0078125,-0.0078125,-0.0078125,-0.0078125,0.0,0.0078125,0.0,-0.015625,-0.046875,0.078125,0.0625,-0.0390625,-0.015625,-0.0390625,0.0078125,-0.0546875,-0.0078125,-0.015625,-0.015625,0.0,0.015625,-0.015625,-0.0546875,-0.0390625,-0.015625,-0.0078125,0.0078125,0.015625,0.0859375,-0.0078125,-0.03125,-0.0234375,-0.0,-0.0234375,-0.0078125,0.0078125,0.0078125,-0.0078125,-0.015625,0.015625,0.0078125,-0.0078125,0.0078125,-0.0390625,0.0078125,-0.0234375,-0.015625,-0.0234375,-0.078125,-0.015625,-0.0546875,-0.0,0.0625,0.109375,-0.0078125,0.0,0.0390625,-0.0546875,-0.0234375,0.0078125,0.0078125,-0.0234375,0.0234375,-0.0078125,0.0,-0.046875,-0.015625,-0.0546875,-0.046875,-0.0078125,0.0078125,0.015625,0.0078125,-0.0,0.0234375,-0.0390625,-0.0078125,0.0390625,-0.0234375,0.0234375,0.0703125,0.0390625,-0.0546875,-0.03125,-0.0390625,0.03125,0.046875,-0.0234375,-0.0,0.03125,-0.0234375,0.015625,0.015625,-0.0234375,-0.015625,0.0078125,-0.0234375,-0.046875,0.0390625,0.0078125,-0.015625,0.015625,0.015625,0.0078125,0.015625,0.0078125,-0.0078125,-0.0,-0.0,-0.0078125,-0.0390625,0.0078125,0.0234375,-0.0390625,0.0078125,-0.0390625,-0.0234375,0.0078125,-0.015625,-0.0234375,0.0234375,-0.015625,0.03125,-0.046875,-0.0546875,-0.0390625,0.0078125,-0.0234375,-0.0546875,0.0546875,0.015625,0.015625,-0.03125,0.0078125,0.0078125,0.0078125,0.0234375,0.015625,0.0078125,0.0,0.0,-0.0,0.0078125,-0.015625,-0.0078125,-0.015625,-0.0,-0.0390625,-0.0078125,0.0,-0.0,-0.0078125,-0.015625,-0.0234375,-0.015625,-0.0234375,0.0078125,0.0703125,-0.0234375,0.0234375,0.015625,0.0078125,0.0,-0.015625,-0.0703125,0.0234375,-0.0390625,-0.0234375,-0.015625,0.0,0.015625,-0.0234375,-0.0625,-0.109375,0.015625,0.109375,0.03125,-0.0078125,-0.015625,0.0234375,-0.0390625,-0.0234375,-0.0078125,0.0,-0.0234375,0.0625,0.0078125,-0.046875,-0.0234375,0.0234375,0.0625,0.0859375,0.0234375,-0.0078125,-0.03125,0.0,-0.015625,0.0078125,-0.03125,-0.015625,-0.03125,0.015625,0.046875,-0.109375,0.078125,-0.0546875,-0.015625,-0.0,-0.0234375,-0.0625,-0.0078125,0.0078125,0.03125,0.0078125,0.0234375,-0.03125,0.03125,0.0546875,-0.0390625,-0.015625,-0.0390625,-0.0078125,0.03125,0.03125,0.0703125,-0.0390625,0.0234375,-0.03125,0.015625,0.0,-0.0390625,0.0234375,-0.0234375,-0.0703125,0.015625,-0.046875,-0.0390625,-0.046875,0.0703125,0.0390625,-0.0546875,0.03125,0.03125,0.046875,0.046875,0.0078125,-0.03125,0.046875,0.0234375,-0.0703125,0.0078125,0.03125,0.0625,-0.015625,0.015625,-0.0234375,-0.03125,-0.03125,0.0234375,0.0078125,-0.015625,0.0078125,0.0390625,-0.0390625,-0.0078125,-0.0390625,-0.0390625,-0.0,0.0078125,0.015625,-0.0390625,-0.03125,0.015625,-0.046875,-0.015625,-0.0078125,0.015625,-0.0546875,-0.0078125,-0.015625,-0.0078125,0.0,0.015625,0.0078125,0.0625,-0.0078125,-0.0078125,0.0078125,-0.0078125,0.0,0.0078125,0.0,0.0,-0.015625,0.0078125,-0.015625,-0.0703125,0.0234375,-0.03125,0.0078125,-0.0234375,-0.0,0.0234375,0.0390625,0.0234375,-0.03125,0.03125,-0.0390625,-0.078125,-0.0078125,0.046875,0.015625,-0.0,0.0078125,0.03125,0.0234375,-0.0703125,0.015625,-0.0546875,0.0390625,-0.0078125,0.0234375,-0.0078125,-0.0078125,-0.015625,-0.0078125,0.0,0.0078125,0.0078125,-0.015625,0.0078125,0.0,-0.0234375,0.03125,-0.015625,0.0,0.0078125,0.0546875,0.015625,0.0234375,-0.078125,-0.0078125,-0.046875,0.0546875,-0.078125,-0.0078125,-0.0078125,-0.03125,0.0703125,-0.0625,0.046875,-0.0234375,-0.0234375,0.015625,-0.0546875,-0.046875,0.09375,-0.0078125,-0.03125,-0.015625,-0.046875,-0.03125,0.0546875,0.015625,-0.0703125,-0.0390625,-0.0390625,0.0390625,0.03125,0.0390625,0.015625,-0.0234375,-0.0390625,-0.046875,0.03125,0.0390625,-0.015625,-0.015625,-0.03125,0.03125,-0.0078125,-0.0390625,0.0546875,0.0078125,0.03125,-0.046875,-0.046875,-0.0078125,0.0390625,0.0078125,-0.015625,0.046875,-0.0078125,0.0,-0.0078125,-0.0078125,0.03125,-0.0234375,-0.0078125,0.03125,-0.0,0.078125,-0.0078125,-0.0078125,0.0390625,0.0078125,-0.03125,-0.1015625,0.03125,0.0546875,-0.03125,0.0703125,0.0390625,-0.0390625,0.0078125,-0.015625,-0.0703125,0.03125,-0.109375,-0.03125,-0.0546875,0.0078125,0.0234375,0.0078125,0.0078125,0.0234375,0.03125,-0.0,0.0,0.0078125,0.015625,0.0078125,-0.0078125,0.015625,0.078125,-0.0078125,0.0078125,0.0546875,0.0078125,0.046875,0.03125,0.0859375,0.0234375,-0.0546875,-0.0234375,0.0625,-0.046875,-0.0078125,0.015625,-0.015625,0.0078125,-0.046875,-0.1015625,-0.0,0.0625,0.09375,0.0390625,-0.0234375,0.015625,0.0390625,0.0234375,-0.0625,-0.046875,0.1015625,0.015625,0.0859375,-0.03125,-0.03125,0.0078125,-0.0234375,-0.0078125,0.0234375,-0.0625,-0.0,-0.0390625,0.015625,-0.03125,0.0390625,-0.015625,0.0625,-0.0703125,0.0546875,0.0078125,-0.0546875,0.03125,-0.0703125,0.0625,0.0625,-0.109375,-0.0078125,0.015625,-0.0546875,0.0234375,-0.0078125,0.09375,0.03125,-0.0546875,0.09375,-0.0,-0.015625,0.0390625,-0.0078125,-0.046875,0.015625,0.0546875,0.0390625,-0.0078125,-0.046875,0.0546875,0.015625,0.046875,-0.03125,-0.0703125,0.03125,0.0234375,-0.0546875,-0.0390625,-0.0703125,-0.03125,-0.0,0.0,-0.0,0.09375,-0.046875,-0.015625,-0.0703125,-0.015625,0.0234375,-0.0234375,0.0390625,0.015625,0.0234375,0.0390625,-0.078125,-0.0390625,0.109375,-0.0703125,0.09375,0.0078125,-0.0625,0.046875,0.03125,-0.0859375,-0.0546875,-0.03125,-0.015625,-0.0390625,-0.015625,-0.0859375,-0.0234375,0.1171875,-0.0625,-0.046875,0.015625,-0.046875,0.0,0.0234375,-0.0234375,0.0234375,0.0234375,-0.0625,-0.03125,-0.0703125,-0.0078125,-0.0,-0.0234375,-0.015625,-0.0,0.0546875,0.046875,0.0234375,-0.09375,-0.0703125,0.015625,0.0078125,-0.0,0.0078125,-0.0078125,0.0,-0.0078125,-0.0078125,-0.015625,-0.0,-0.015625,-0.015625,-0.0390625,0.046875,-0.0234375,-0.0234375,0.0625,0.0,-0.0078125,-0.0390625,0.015625,0.0078125,0.046875,-0.0234375,0.046875,0.046875,-0.015625,0.0078125,0.0234375,0.0546875,0.03125,0.0078125,-0.0703125,0.015625,-0.015625,-0.0078125,-0.03125,-0.0078125,-0.0078125,-0.0078125,-0.0078125,-0.0,0.0078125,-0.015625,-0.0078125,0.0078125,-0.0234375,-0.0078125,-0.015625,0.0390625,0.0234375,0.0546875,0.046875,-0.015625,-0.0078125,-0.0078125,0.078125,0.0546875,-0.0390625,-0.0,0.0390625,-0.015625,0.0078125,-0.0078125,-0.0078125,0.046875,0.015625,-0.046875,-0.015625,-0.0390625,0.0390625,-0.015625,-0.0234375,0.015625,-0.0390625,-0.0625,0.0078125,0.015625,-0.0234375,-0.046875,-0.0546875,-0.03125,-0.0078125,0.0078125,0.015625,0.078125,-0.03125,0.046875,-0.078125,-0.0078125,0.015625,0.015625,-0.0,0.0234375,-0.046875,0.0703125,0.015625,-0.0078125,0.0078125,0.015625,0.0078125,-0.0,-0.0,-0.03125,0.03125,-0.03125,0.0078125,0.0,0.0078125,-0.0234375,0.0390625,-0.0234375,-0.078125,-0.03125,-0.0234375,0.0078125,0.03125,0.015625,-0.0546875,-0.0234375,-0.046875,0.0859375,0.0546875,0.0078125,-0.0390625,-0.0625,0.0078125,0.015625,-0.0234375,-0.015625,0.1328125,-0.015625,-0.09375,0.0625,-0.0078125,0.0078125,-0.0,-0.0,0.015625,0.03125,-0.015625,0.015625,0.0234375,-0.0078125,0.0,-0.0390625,-0.015625,-0.0234375,0.0078125,-0.015625,0.0234375,0.0234375,0.0078125,-0.015625,-0.03125,-0.0078125,-0.015625,0.0546875,0.0,-0.03125,0.0234375,-0.0078125,-0.046875,0.015625,-0.0234375,-0.03125,-0.0546875,0.03125,-0.03125,0.0234375,0.015625,-0.015625,-0.0390625,-0.046875,-0.015625,0.03125,-0.0234375,-0.0234375,0.0703125,0.078125,0.03125,0.046875,-0.046875,0.0,-0.0234375,0.03125,-0.0078125,0.015625,-0.046875,-0.046875,0.0078125,-0.0,-0.0078125,0.1328125,-0.0234375,0.0546875,0.09375,0.0,-0.0,-0.0234375,-0.0,0.015625,-0.0390625,-0.0625,-0.0625,0.1328125,0.0859375,-0.046875,-0.0390625,-0.0625,0.03125,-0.0625,-0.0703125,-0.0234375,0.0078125,0.015625,0.0078125,0.078125,0.078125,0.015625,-0.0234375,0.0234375,0.015625,-0.0078125,-0.0390625,-0.0390625,0.046875,-0.0,0.015625,-0.0078125,0.109375,-0.0546875,-0.0,-0.0078125,-0.015625,-0.0234375,0.078125,0.0234375,-0.109375,-0.015625,-0.0390625,0.0546875,-0.015625,-0.0078125,-0.0078125,0.0546875,-0.0390625,-0.0078125,-0.0625,-0.046875,-0.0546875,-0.0390625,-0.03125,0.078125,-0.0234375,0.0,0.0078125,-0.0703125,0.015625,0.015625,0.0078125,-0.046875,0.046875,-0.0625,-0.0546875,-0.0,-0.0234375,-0.03125,0.0078125,0.015625,0.0078125,-0.0625,-0.0234375,0.015625,-0.0625,-0.0625,-0.015625,0.0078125,0.0,-0.0390625,0.0,0.0390625,0.0703125,-0.015625,0.0703125,-0.03125,-0.015625,-0.0078125,-0.0703125,0.0078125,-0.0,-0.0078125,0.0078125,0.015625,0.0078125,0.015625,0.0,0.015625,-0.0,-0.0,-0.0234375,-0.03125,-0.109375,-0.09375,0.0234375,0.015625,0.109375,-0.03125,0.03125,-0.0,-0.0546875,-0.0390625,0.0078125,-0.0546875,0.046875,0.0234375,0.015625,-0.0,0.0078125,-0.015625,0.0234375,-0.0703125,-0.0390625,-0.0078125,0.0234375,-0.0078125,0.0,-0.0078125,0.0078125,-0.0078125,0.0234375,0.0,0.0078125,-0.0078125,-0.0,-0.0546875,-0.0234375,-0.0703125,-0.0234375,-0.0546875,-0.015625,0.15625,-0.0390625,0.0,0.0234375,-0.0703125,-0.0078125,-0.1796875,0.15625,-0.0078125,-0.1015625,0.0546875,0.0078125,-0.0234375,0.0625,0.0078125,0.0234375,0.03125,-0.0625,0.0234375,-0.0859375,0.015625,0.015625,-0.0078125,-0.0078125,-0.0859375,0.0390625,0.0078125,-0.015625,-0.0234375,-0.015625,-0.0546875,0.0234375,-0.0234375,0.0859375,0.046875,0.03125,0.1171875,-0.078125,0.015625,0.0,-0.03125,-0.03125,0.0078125,0.0078125,0.015625,-0.03125,-0.0,-0.0234375,0.0234375,0.046875,0.0078125,-0.03125,0.0,-0.0078125,-0.0234375,-0.0078125,0.015625,0.0078125,-0.046875,0.0078125,-0.0234375,0.0,0.0234375,0.046875,0.0859375,-0.0078125,-0.03125,0.0234375,-0.0546875,0.0078125,-0.09375,-0.015625,0.0234375,0.0859375,-0.0234375,-0.0,0.1015625,-0.0234375,-0.03125,-0.0234375,-0.046875,-0.015625,-0.1015625,-0.0078125,0.0078125,-0.0,-0.0078125,-0.0,-0.0,0.0,-0.0078125,-0.03125,-0.0078125,0.0234375,-0.0390625,0.0078125,-0.0078125,-0.0078125,0.0078125,0.0,0.03125,-0.0078125,0.0390625,-0.03125,-0.0234375,0.046875,0.03125,-0.0703125,0.0078125,-0.0078125,-0.0078125,-0.078125,-0.078125,-0.046875,0.0390625,0.0234375,-0.03125,-0.09375,0.2109375,0.0390625,0.0703125,0.0546875,0.0,-0.0078125,-0.0703125,-0.015625,-0.0078125,0.046875,-0.03125,0.015625,0.015625,-0.0390625,-0.046875,-0.0859375,0.015625,0.03125,-0.0390625,-0.0078125,0.03125,0.0703125,-0.0390625,0.0078125,-0.0546875,-0.03125,-0.03125,-0.015625,-0.0390625,0.0703125,-0.1015625,-0.046875,0.0390625,0.0234375,-0.0234375,-0.09375,0.109375,0.0078125,-0.03125,0.0078125,-0.0078125,0.0546875,0.0625,-0.03125,0.015625,-0.046875,-0.0234375,-0.0078125,0.0234375,0.015625,-0.03125,-0.0078125,-0.015625,-0.0234375,-0.015625,-0.0546875,-0.0625,-0.1171875,-0.0625,-0.03125,0.0625,-0.0234375,0.0078125,0.0625,0.0625,0.0546875,-0.015625,-0.0234375,-0.109375,-0.03125,-0.0234375,0.0546875,-0.0234375,0.0234375,0.078125,-0.0234375,-0.0390625,-0.03125,-0.0234375,-0.03125,0.015625,0.0703125,-0.0234375,-0.046875,-0.0078125,0.015625,-0.03125,-0.03125,0.0390625,-0.0625,0.03125,-0.0078125,0.03125,0.0546875,0.0,-0.0,-0.0,-0.03125,-0.0234375,0.046875,-0.0,-0.015625,-0.078125,-0.015625,-0.046875,0.09375,-0.03125,-0.046875,0.0234375,-0.0390625,-0.015625,-0.0234375,0.015625,-0.015625,-0.03125,0.046875,-0.0234375,0.03125,-0.015625,-0.015625,-0.015625,-0.015625,-0.015625,-0.0078125,0.015625,0.0078125,0.0078125,-0.015625,0.0078125,-0.046875,-0.0234375,-0.0546875,0.0,0.078125,0.046875,-0.015625,0.015625,0.015625,-0.046875,0.0078125,-0.015625,0.015625,0.015625,0.0859375,-0.0078125,-0.0234375,-0.0078125,-0.0,-0.0,-0.0546875,0.0078125,0.078125,-0.0546875,0.09375,0.0,0.0078125,0.0078125,-0.0078125,-0.0,0.0078125,0.0,0.0078125,0.0,-0.0078125,0.015625,0.03125,-0.0390625,-0.0546875,0.0234375,-0.0390625,0.1328125,-0.046875,-0.0546875,0.03125,-0.03125,-0.09375,0.0859375,0.0078125,-0.0546875,0.03125,0.09375,0.078125,-0.03125,0.0078125,0.0859375,-0.109375,-0.0078125,0.0234375,0.0,-0.0546875,0.0546875,-0.0234375,0.0234375,-0.0390625,0.015625,-0.0234375,0.0078125,0.0234375,-0.0234375,0.03125,-0.0234375,-0.015625,0.0234375,-0.0546875,0.015625,-0.0234375,-0.015625,0.0078125,-0.015625,-0.015625,0.03125,-0.015625,0.03125,-0.0390625,0.0,-0.0078125,0.03125,-0.03125,-0.046875,0.015625,0.0078125,-0.0,0.0078125,0.015625,-0.0078125,-0.015625,0.0546875,0.046875,-0.0078125,0.0234375,-0.0,-0.0234375,0.015625,-0.0078125,-0.015625,0.015625,0.0078125,0.015625,0.0390625,-0.0625,-0.0390625,-0.0078125,0.09375,0.0078125,-0.015625,-0.0078125,-0.0078125,0.0390625,-0.03125,-0.078125,0.0078125,0.015625,-0.046875,-0.0078125,-0.0,-0.0078125,-0.0078125,-0.0078125,0.015625,-0.0078125,-0.0078125,-0.015625,0.015625,0.015625,0.015625,-0.0078125,0.015625,0.015625,-0.0234375,0.0625,-0.0,0.0390625,0.0078125,0.0,-0.0234375,-0.0234375,0.0,-0.03125,-0.046875,0.03125,-0.03125,-0.0,0.0078125,-0.015625,-0.0546875,-0.0078125,-0.0078125,-0.015625,-0.046875,0.0078125,-0.0546875,-0.046875,-0.03125,-0.0625,0.0078125,-0.046875,-0.0859375,0.046875,-0.015625,-0.0234375,0.0625,-0.0078125,0.03125,-0.03125,0.0703125,-0.078125,0.0234375,0.015625,0.046875,-0.03125,0.03125,-0.0390625,-0.0078125,-0.0078125,0.046875,-0.015625,0.1015625,0.0,-0.0078125,-0.046875,-0.03125,0.015625,0.0234375,-0.03125,0.0234375,0.015625,0.0390625,0.0546875,-0.0390625,-0.0078125,-0.0078125,0.015625,0.03125,0.0390625,0.0546875,0.0234375,-0.0078125,0.03125,-0.0390625,0.0234375,-0.0234375,-0.015625,0.0390625,0.0234375,-0.03125,-0.0390625,0.0390625,0.0234375,-0.0234375,0.0,-0.03125,-0.0234375,0.109375,0.0234375,0.0390625,-0.0234375,-0.0546875,-0.0390625,-0.0625,-0.015625,-0.015625,0.0234375,-0.0234375,-0.03125,-0.0703125,-0.015625,-0.046875,0.0390625,-0.0078125,0.0546875,-0.015625,0.015625,-0.0546875,0.046875,0.0078125,0.0,0.015625,0.0546875,0.0390625,-0.0546875,0.0078125,-0.078125,-0.03125,-0.0625,-0.0,-0.0078125,0.046875,0.0078125,0.015625,0.046875,-0.015625,0.0078125,-0.046875,0.0,-0.0,-0.0234375,0.0859375,0.0234375,0.0,0.0,-0.046875,-0.046875,-0.0234375,-0.0,-0.0078125,-0.015625,0.0078125,-0.0078125,0.0078125,0.0078125,-0.015625,-0.015625,-0.015625,-0.0078125,0.015625,-0.046875,-0.0234375,-0.046875,0.0390625,0.0390625,-0.0234375,-0.0625,-0.046875,-0.0078125,0.0390625,0.015625,-0.0078125,-0.0078125,-0.0078125,-0.015625,-0.0625,-0.0625,-0.015625,0.0234375,0.078125,-0.0,0.0078125,0.0078125,0.0078125,-0.0078125,-0.046875,0.0234375,-0.0078125,0.0078125,-0.0078125,0.0078125,0.0078125,0.0,-0.0078125,-0.0078125,-0.0,0.09375,0.015625,-0.0234375,-0.0390625,-0.015625,0.0078125,-0.0546875,-0.078125,-0.046875,-0.0234375,-0.0078125,0.03125,0.1953125,0.0703125,-0.03125,0.0625,0.0078125,0.03125,0.0234375,-0.0390625,-0.0078125,0.1171875,0.0625,0.0078125,-0.015625,-0.0625,-0.046875,-0.0078125,-0.0234375,-0.0,0.015625,-0.015625,0.0078125,0.0078125,-0.0390625,0.015625,-0.015625,-0.046875,-0.0078125,-0.0234375,-0.0546875,-0.015625,0.0546875,-0.0,-0.0234375,0.0546875,0.0078125,0.015625,0.015625,0.015625,-0.0078125,-0.0,-0.03125,-0.015625,-0.03125,-0.0078125,-0.0,0.0234375,0.0703125,0.0078125,-0.015625,0.0,0.0234375,0.0234375,0.0390625,0.0078125,-0.046875,0.015625,0.015625,-0.0390625,-0.0390625,-0.03125,-0.1015625,-0.1171875,-0.0078125,-0.0390625,-0.0390625,-0.0234375,0.0234375,-0.0078125,-0.0078125,0.0390625,0.0234375,-0.046875,0.0234375,-0.0078125,-0.015625,-0.03125,0.03125,0.0625,-0.015625,0.0,0.015625,0.0078125,-0.015625,-0.0,0.0,-0.015625,0.0078125,0.015625,0.0,-0.0078125,-0.0078125,-0.0546875,0.0078125,0.0234375,-0.0,-0.0234375,-0.015625,-0.0234375,-0.015625,0.0,0.0,-0.03125,-0.0078125,-0.0078125,0.046875,0.0546875,-0.0078125,-0.0234375,-0.0,-0.0234375,-0.015625,-0.0546875,-0.078125,0.03125,0.0078125,0.0,-0.0,-0.0,-0.0234375,-0.015625,-0.0234375,0.046875,0.015625,0.0,-0.0390625,0.015625,-0.0625,-0.03125,-0.03125,-0.0859375,-0.0625,0.0234375,-0.03125,-0.0,-0.0234375,0.046875,0.015625,-0.0390625,-0.015625,0.046875,-0.015625,-0.015625,-0.0234375,-0.0234375,-0.0625,0.0078125,-0.0078125,-0.0390625,-0.0,0.0546875,-0.0546875,-0.0234375,-0.0078125,-0.0703125,-0.078125,-0.0234375,0.0390625,0.015625,-0.0625,-0.0234375,-0.015625,0.0,-0.0390625,0.0625,0.0625,-0.0078125,-0.0625,0.0078125,0.0703125,0.0625,0.0234375,-0.078125,-0.0625,0.0234375,-0.0390625,0.0078125,0.0078125,-0.0546875,0.0078125,-0.046875,0.0859375,0.03125,0.03125,0.046875,-0.0078125,-0.046875,-0.015625,-0.046875,-0.0234375,0.0078125,-0.0859375,-0.0234375,-0.0625,0.0234375,0.0,-0.03125,-0.0234375,-0.0078125,-0.0078125,0.0,0.0390625,-0.0,-0.015625,-0.0234375,-0.046875,-0.0234375,0.0234375,0.0703125,-0.0078125,-0.046875,0.0390625,0.1171875,0.0390625,-0.0390625,-0.0390625,0.0,0.03125,-0.0234375,-0.015625,0.109375,-0.0625,0.015625,-0.03125,0.0078125,-0.0,-0.0,-0.0234375,-0.046875,-0.0234375,-0.0625,-0.0859375,0.0,-0.0078125,0.0078125,0.0078125,0.0,0.015625,0.0078125,-0.015625,-0.0078125,-0.0078125,0.03125,0.0390625,0.09375,-0.09375,-0.015625,-0.0859375,0.03125,-0.015625,-0.015625,0.015625,0.0078125,0.046875,-0.0703125,-0.046875,-0.03125,-0.0390625,0.078125,-0.03125,-0.015625,0.0078125,-0.09375,-0.03125,0.0859375,-0.0703125,0.0859375,0.140625,-0.0,0.0078125,-0.0078125,-0.0,0.0078125,-0.0,-0.0,0.0078125,0.0,0.09375,-0.0546875,0.0859375,-0.0234375,0.015625,-0.1328125,-0.03125,0.1328125,-0.09375,-0.0390625,-0.0390625,-0.1015625,-0.03125,0.0,0.0234375,-0.0390625,-0.03125,0.1328125,0.0,-0.078125,-0.078125,0.015625,0.125,-0.078125,-0.0859375,-0.0234375,0.0390625,0.03125,-0.0234375,-0.0390625,0.0625,-0.09375,-0.0234375,0.0390625,-0.0078125,-0.015625,0.03125,-0.0546875,-0.0390625,-0.0390625,0.03125,-0.078125,-0.0078125,0.109375,0.1015625,-0.0078125,0.0078125,0.0390625,0.0,0.078125,0.09375,0.0390625,-0.0234375,-0.0625,0.0234375,0.03125,-0.015625,0.046875,0.0234375,-0.0234375,-0.0078125,0.0546875,-0.015625,0.0078125,-0.015625,0.015625,-0.046875,-0.0703125,-0.03125,-0.0625,0.0390625,-0.0703125,-0.0234375,-0.0546875,0.03125,-0.0078125,0.046875,0.0390625,-0.0703125,-0.0390625,0.0390625,-0.015625,-0.0234375,0.0859375,-0.03125,-0.109375,0.0390625,0.046875,-0.109375,-0.0078125,-0.0078125,0.0078125,0.015625,-0.015625,-0.0234375,0.0,-0.0078125,-0.0078125,0.0,-0.03125,-0.0078125,0.015625,0.0703125,-0.0859375,-0.015625,0.03125,-0.0390625,-0.046875,-0.03125,0.0234375,-0.0234375,0.0078125,-0.046875,0.015625,0.0078125,-0.0625,-0.0234375,0.015625,-0.0546875,-0.078125,0.0390625,0.0234375,0.015625,0.0,-0.015625,-0.015625,-0.015625,-0.0859375,-0.09375,0.0078125,-0.0,0.0859375,0.015625,-0.0078125,0.0078125,0.0234375,-0.015625,0.0234375,0.015625,-0.03125,0.0859375,-0.0,-0.0546875,-0.0546875,-0.015625,0.03125,0.015625,0.0078125,-0.0625,0.03125,0.0234375,0.0078125,-0.0546875,-0.078125,-0.0,0.0546875,0.0703125,0.0078125,0.0546875,0.0234375,-0.03125,-0.0703125,-0.015625,0.0078125,0.0,-0.0078125,0.0859375,0.015625,-0.0,0.0078125,0.0546875,0.0,0.0078125,-0.046875,-0.109375,0.015625,-0.0078125,-0.0390625,0.078125,0.078125,0.0546875,-0.015625,-0.0703125,0.09375,-0.0078125,-0.0703125,0.078125,-0.015625,-0.0546875,-0.1015625,-0.078125,0.03125,0.015625,-0.0390625,0.0703125,-0.015625,0.0703125,-0.1875,-0.03125,-0.03125,-0.015625,-0.0546875,-0.0078125,-0.015625,-0.1171875,0.0078125,-0.0234375,-0.0,0.0,0.0078125,0.0234375,-0.0625,-0.09375,-0.0078125,-0.0,-0.015625,-0.0234375,-0.0546875,-0.078125,0.0703125,-0.015625,-0.0078125,0.0078125,-0.015625,-0.015625,-0.1015625,-0.09375,-0.015625,0.0625,0.015625,-0.0078125,0.1796875,-0.0859375,-0.0234375,-0.015625,0.0703125,-0.0,-0.0390625,-0.0,-0.0859375,-0.015625,-0.0078125,-0.046875,0.0078125,0.0,-0.0078125,-0.0078125,0.0078125,-0.0078125,0.0,0.0078125,-0.015625,0.0390625,0.0390625,0.0078125,-0.0,0.0234375,0.0078125,-0.0546875,-0.0625,-0.078125,0.0,0.03125,-0.015625,-0.0,0.0078125,0.015625,0.0078125,0.0078125,-0.0078125,-0.015625,0.015625,-0.046875,-0.03125,0.0078125,0.03125,0.1015625,0.0234375,-0.015625,-0.0078125,-0.0078125,-0.0,0.0,0.0078125,0.0078125,-0.0078125,-0.015625,-0.0078125,-0.015625,0.0,-0.0078125,-0.0390625,-0.0234375,-0.03125,-0.0234375,0.046875,-0.0390625,-0.0546875,-0.078125,0.0625,0.015625,-0.0546875,-0.078125,0.1015625,-0.09375,-0.0390625,0.015625,0.0390625,0.078125,0.0,-0.078125,0.03125,-0.03125,0.0234375,0.03125,0.0234375,0.0078125,0.0078125,0.03125,0.046875,-0.015625,-0.0078125,-0.046875,-0.046875,-0.0078125,0.0234375,0.0390625,-0.046875,-0.0234375,-0.0546875,0.0234375,0.125,-0.0078125,-0.0078125,0.0078125,0.0078125,0.015625,0.0546875,-0.0390625,-0.0390625,-0.03125,0.0,0.015625,-0.03125,0.0234375,0.0078125,-0.0234375,0.0,0.0234375,0.0078125,0.015625,0.0,-0.0234375,0.0078125,-0.0234375,-0.03125,0.09375,-0.03125,0.0390625,0.015625,0.0078125,-0.046875,-0.03125,-0.0546875,0.09375,0.0390625,-0.0234375,-0.0625,0.0078125,0.03125,-0.0703125,0.0078125,-0.0390625,0.03125,-0.1015625,-0.0546875,0.0703125,-0.0,0.015625,0.0078125,0.0,0.0078125,-0.015625,-0.015625,-0.0078125,-0.0078125,0.0,-0.0078125,0.046875,-0.0078125,-0.015625,-0.0390625,-0.03125,-0.0078125,-0.0234375,0.0078125,-0.0390625,-0.0625,-0.046875,-0.015625,0.1171875,-0.0078125,0.0078125,-0.0078125,-0.0703125,-0.03125,-0.046875,0.015625,-0.046875,-0.0234375,0.0078125,-0.046875,0.0,-0.0078125,-0.03125,0.0078125,-0.0390625,-0.0390625,0.0234375,0.015625,-0.03125,0.046875,0.015625,0.046875,-0.015625,-0.046875,0.0390625,0.0234375,-0.03125,-0.0078125,-0.03125,-0.078125,0.015625,-0.0234375,-0.1015625,0.015625,-0.03125,0.0,0.0,-0.046875,-0.0703125,-0.0390625,-0.0625,-0.015625,-0.03125,-0.046875,0.1015625,-0.0234375,-0.015625,-0.046875,-0.015625,0.0,0.0078125,-0.0390625,-0.015625,-0.0703125,0.03125,0.0234375,-0.0703125,-0.0078125,-0.03125,-0.0625,0.0234375,0.046875,-0.0234375,0.0390625,-0.015625,-0.0078125,0.015625,-0.03125,0.0390625,-0.015625,-0.0234375,0.0625,-0.0390625,-0.0546875,-0.0234375,-0.0078125,-0.0,-0.0546875,-0.0,0.046875,0.078125,0.03125,0.0078125,0.0546875,-0.0546875,-0.09375,-0.0390625,-0.015625,-0.015625,0.109375,0.0078125,-0.0,-0.0390625,-0.015625,0.0,0.0390625,0.0078125,-0.03125,-0.046875,0.015625,0.015625,-0.046875,-0.03125,-0.0234375,-0.046875,0.03125,-0.0390625,-0.03125,-0.0078125,0.015625,-0.015625,-0.03125,-0.015625,0.078125,0.0078125,0.015625,-0.046875,-0.0,-0.0234375,-0.0078125,-0.0625,0.0859375,0.03125,-0.03125,-0.03125,-0.0234375,0.0234375,-0.0546875,-0.09375,-0.0,-0.0078125,-0.0078125,-0.0078125,0.0078125,-0.015625,-0.015625,-0.0,0.0078125,-0.0,0.046875,0.109375,-0.0078125,-0.0546875,0.0234375,-0.046875,0.0234375,0.03125,-0.03125,-0.0234375,0.0,-0.0546875,-0.0703125,0.0546875,-0.015625,0.0078125,0.0859375,0.0234375,-0.0859375,0.0078125,0.015625,-0.078125,-0.015625,-0.0390625,0.171875,-0.0390625,0.0078125,-0.0078125,-0.015625,0.0078125,0.0,-0.0078125,0.0078125,0.0,0.0078125,-0.046875,-0.046875,-0.0859375,-0.1015625,-0.046875,0.03125,0.03125,-0.0078125,0.03125,0.09375,-0.0234375,-0.03125,-0.0390625,-0.0078125,-0.0078125,-0.0234375,0.0,-0.0546875,0.0,-0.0078125,0.0,-0.0078125,0.015625,0.0859375,-0.0078125,0.0546875,-0.1015625,-0.046875,-0.03125,0.078125,0.03125,-0.015625,-0.0234375,-0.0,-0.0234375,-0.015625,0.015625,-0.015625,-0.0625,-0.0546875,-0.015625,0.078125,-0.0703125,-0.0546875,-0.0390625,-0.0078125,-0.03125,-0.015625,-0.0078125,-0.0,0.0078125,-0.015625,-0.03125,-0.0546875,0.015625,-0.0078125,-0.015625,-0.0234375,0.0078125,0.0078125,0.046875,0.03125,0.0078125,0.0078125,-0.015625,-0.0625,-0.0078125,0.0234375,0.046875,-0.046875,0.0078125,-0.015625,-0.0078125,0.0625,0.046875,-0.015625,-0.0390625,0.0234375,0.015625,-0.15625,-0.046875,-0.0234375,-0.0234375,0.0703125,0.0390625,-0.015625,-0.03125,0.015625,0.0234375,0.03125,-0.0,0.0078125,0.0,-0.015625,-0.015625,-0.0,-0.0078125,0.015625,0.0078125,0.0,-0.0546875,-0.0078125,0.0234375,-0.0546875,-0.0390625,-0.0390625,0.046875,-0.0078125,0.0078125,-0.0078125,-0.0390625,0.03125,0.0625,0.0625,-0.015625,-0.046875,0.0546875,0.03125,0.0,0.03125,-0.03125,0.015625,0.0234375,0.0546875,-0.0234375,-0.0234375,0.0078125,-0.03125,0.0,0.0390625,-0.015625,0.046875,-0.1015625,-0.0625,0.015625,-0.046875,-0.03125,0.0234375,-0.0078125,0.015625,0.046875,-0.0234375,0.0078125,0.0234375,-0.03125,0.0078125,-0.0234375,-0.0625,0.0,-0.015625,-0.0234375,0.015625,-0.0,0.046875,-0.0703125,-0.0703125,-0.0390625,0.0703125,0.0078125,0.0,-0.015625,0.0234375,-0.0078125,-0.0234375,-0.015625,0.03125,-0.078125,-0.015625,-0.0078125,0.0234375,-0.0078125,0.0234375,0.0390625,0.0546875,-0.046875,-0.0546875,-0.0078125,-0.015625,0.046875,-0.0546875,0.0546875,0.0390625,-0.046875,0.0078125,-0.0546875,0.046875,0.0,0.0390625,-0.0234375,-0.0078125,-0.0234375,-0.0,0.0546875,0.109375,0.0078125,-0.0078125,-0.046875,-0.0078125,-0.0,-0.0390625,0.0234375,-0.0546875,-0.0234375,0.0078125,-0.046875,0.015625,-0.046875,0.03125,-0.0078125,-0.03125,-0.0859375,-0.0703125,0.015625,-0.0234375,-0.015625,0.0859375,0.0625,0.0078125,-0.0703125,0.0,-0.046875,0.0078125,0.0390625,-0.0234375,0.03125,0.0234375,-0.0234375,0.0234375,0.0390625,0.0,-0.0,0.0,0.0234375,0.0859375,-0.03125,-0.03125,0.0,0.125,-0.0390625,-0.0,-0.0546875,-0.0625,0.015625,0.0,-0.0078125,-0.015625,-0.0078125,0.0234375,0.0078125,0.0078125,0.0078125,0.0078125,0.0390625,-0.0234375,0.015625,-0.0,0.03125,0.0234375,-0.015625,-0.0625,0.03125,-0.0234375,-0.0625,-0.03125,0.1171875,-0.0234375,-0.015625,0.0546875,-0.0078125,0.0859375,-0.03125,0.078125,0.0234375,0.0234375,-0.03125,-0.015625,0.078125,0.0546875,0.0625,0.0,-0.0078125,0.0078125,-0.015625,-0.0078125,-0.0078125,-0.0078125,0.0,-0.0,0.0390625,0.0546875,-0.0078125,0.1171875,-0.0078125,-0.0546875,-0.109375,0.0703125,0.046875,0.0078125,-0.046875,-0.0078125,-0.0078125,0.015625,-0.0390625,-0.0390625,-0.015625,0.0625,0.078125,0.0078125,-0.03125,0.0,-0.0078125,-0.078125,-0.0546875,-0.046875,0.078125,0.0078125,-0.046875,0.0078125,0.0390625,0.015625,0.0078125,0.0078125,-0.078125,-0.03125,0.0,-0.0078125,-0.015625,-0.046875,-0.0546875,-0.0078125,0.0859375,-0.03125,-0.015625,0.0234375,0.015625,-0.0078125,-0.0546875,-0.0,-0.0078125,-0.015625,-0.0234375,-0.03125,0.03125,-0.015625,-0.015625,0.03125,-0.015625,-0.015625,-0.0390625,0.015625,-0.015625,-0.0234375,-0.0,0.0234375,-0.0546875,0.03125,-0.015625,0.046875,-0.0234375,-0.015625,-0.0234375,0.0078125,-0.015625,0.0546875,-0.046875,-0.0859375,0.0390625,-0.0625,-0.03125,-0.0234375,0.0234375,-0.0625,-0.078125,0.015625,-0.0,0.0859375,-0.0390625,0.0078125,0.0078125,0.0078125,-0.0,-0.0,-0.0078125,-0.0234375,0.0078125,-0.0078125,0.0078125,-0.0234375,0.0390625,0.0078125,0.0,-0.015625,0.0234375,0.0078125,0.0078125,0.0078125,-0.03125,-0.03125,-0.0078125,0.125,-0.078125,0.0390625,-0.0390625,-0.0234375,-0.015625,0.0078125,-0.03125,0.0078125,-0.03125,0.0234375,-0.0234375,-0.015625,0.0390625,-0.0546875,0.03125,-0.03125,-0.03125,-0.078125,-0.0703125,-0.015625,0.078125,0.03125,-0.078125,-0.03125,-0.015625,-0.015625,-0.0625,-0.078125,0.03125,0.0703125,0.0625,-0.0,-0.015625,0.015625,-0.0,0.0703125,-0.0390625,-0.015625,-0.0703125,-0.046875,-0.046875,-0.0625,-0.09375,0.015625,-0.03125,-0.0625,0.03125,0.1171875,0.0390625,-0.0625,0.0546875,0.0078125,-0.0078125,0.015625,0.0078125,-0.0390625,-0.0,0.0078125,0.0078125,-0.046875,-0.0625,-0.03125,-0.03125,-0.0234375,0.046875,0.0,-0.0703125,0.046875,0.015625,-0.0390625,-0.015625,0.0,0.0234375,-0.03125,-0.0859375,0.046875,-0.03125,0.0,0.0625,0.0234375,0.015625,-0.03125,-0.078125,0.125,-0.0703125,-0.0078125,-0.0859375,0.0078125,-0.0078125,0.046875,0.046875,-0.09375,0.0625,0.125,-0.0390625,-0.046875,-0.0234375,-0.03125,-0.0,-0.03125,-0.0546875,0.0390625,-0.078125,-0.015625,-0.015625,-0.0234375,-0.03125,0.0859375,-0.015625,-0.046875,-0.0859375,-0.0546875,0.0625,-0.0625,-0.0234375,-0.015625,0.0234375,-0.03125,-0.015625,0.046875,-0.0234375,-0.0546875,-0.0390625,0.0625,-0.078125,-0.0546875,0.0234375,-0.0078125,-0.0390625,0.0078125,-0.046875,-0.0078125,0.0,0.0,0.0078125,0.0,0.0,0.0,-0.0078125,-0.015625,-0.0078125,-0.015625,0.0078125,0.0078125,-0.0859375,0.0546875,-0.0390625,-0.078125,0.0625,-0.03125,-0.078125,0.078125,0.03125,0.0,-0.1171875,-0.0546875,-0.03125,0.0859375,-0.015625,0.015625,-0.0078125,-0.03125,-0.0859375,0.0390625,-0.0234375,-0.09375,0.0390625,-0.015625,0.0078125,-0.0,-0.0078125,0.0,0.0078125,0.0078125,0.0,-0.015625,0.0546875,-0.0,0.046875,-0.03125,0.0546875,-0.09375,-0.03125,-0.0234375,-0.0625,0.0625,-0.015625,-0.1015625,0.03125,-0.078125,0.0703125,-0.0703125,-0.015625,0.0,-0.0234375,-0.015625,-0.0703125,-0.0546875,0.0390625,0.046875,-0.0234375,-0.0546875,0.109375,-0.03125,0.0234375,-0.03125,0.0,-0.046875,-0.0078125,0.0078125,0.046875,-0.0234375,-0.0234375,0.046875,0.046875,-0.0390625,0.046875,-0.015625,-0.046875,0.03125,0.015625,-0.015625,-0.0078125,-0.0546875,0.015625,0.0703125,0.0234375,0.0078125,-0.0234375,0.0,0.015625,-0.0078125,-0.0078125,0.015625,0.0546875,0.015625,0.0078125,-0.015625,-0.046875,0.015625,-0.0390625,0.0859375,-0.03125,-0.078125,0.046875,0.046875,-0.046875,-0.0,-0.0078125,0.015625,-0.0625,-0.0703125,0.03125,0.0234375,0.0390625,-0.015625,0.015625,-0.0390625,0.1015625,0.0234375,-0.0234375,-0.0703125,0.1015625,0.0625,-0.03125,-0.0078125,-0.015625,-0.03125,-0.015625,-0.015625,0.0,0.0234375,-0.0078125,0.015625,0.0390625,0.0,-0.0234375,-0.0390625,0.0078125,-0.0078125,-0.015625,-0.0078125,0.03125,0.03125,-0.078125,-0.015625,0.0078125,0.015625,-0.046875,-0.015625,-0.03125,-0.0234375,-0.015625,0.0546875,0.0234375,-0.0546875,0.0078125,-0.0546875,0.0625,0.0234375,0.03125,0.0234375,-0.0078125,0.0390625,-0.0390625,0.0078125,-0.046875,-0.0078125,0.03125,0.0859375,-0.0390625,-0.0078125,-0.0078125,-0.0703125,-0.015625,-0.0,-0.0625,-0.0390625,0.0234375,0.0234375,-0.0390625,-0.0625,-0.09375,-0.0390625,-0.0546875,0.0234375,-0.0234375,0.0390625,0.078125,0.0390625,-0.0703125,0.046875,0.0234375,-0.09375,0.09375,-0.0234375,0.0078125,0.140625,-0.03125,0.03125,-0.0703125,0.0,-0.0703125,0.0234375,0.0,0.0,0.015625,-0.0078125,-0.0,0.03125,-0.0625,-0.0390625,0.1171875,0.0,-0.0078125,0.0078125,0.0703125,-0.0546875,0.0078125,0.0390625,0.0234375,0.0078125,-0.0625,-0.015625,0.1484375,-0.078125,0.0234375,0.1328125,-0.0390625,-0.1640625,0.109375,0.1171875,0.03125,-0.0703125,-0.0390625,0.0234375,0.0234375,-0.015625,0.0234375,-0.046875,-0.0546875,-0.0078125,-0.0390625,-0.015625,-0.109375,0.09375,0.0703125,-0.0859375,-0.03125,-0.0546875,-0.0390625,0.03125,-0.015625,-0.0546875,-0.0625,0.0546875,-0.09375,0.0625,-0.046875,-0.0546875,0.0234375,-0.0078125,0.046875,-0.0,-0.03125,0.03125,-0.03125,-0.1015625,-0.0390625,-0.0546875,0.0078125,0.0078125,-0.0234375,-0.015625,0.03125,0.0,-0.0390625,-0.0078125,0.015625,0.0078125,0.0078125,-0.0078125,-0.0078125,-0.015625,-0.0,-0.0,0.0078125,-0.0078125,0.0234375,-0.0234375,-0.0078125,0.046875,0.015625,0.015625,-0.0078125,-0.0234375,-0.0390625,0.0,0.03125,-0.03125,0.03125,-0.03125,0.03125,0.0234375,-0.03125,-0.0234375,0.0390625,0.03125,0.03125,0.0390625,-0.0078125,-0.0078125,-0.0234375,-0.0078125,-0.0078125,-0.0,0.0,0.0078125,-0.015625,-0.0,-0.0078125,-0.0,0.0078125,-0.0078125,0.0234375,0.0234375,0.015625,0.0390625,-0.0390625,-0.0234375,-0.0390625,-0.046875,0.0625,-0.015625,0.0,0.0234375,0.015625,-0.0078125,-0.015625,0.0390625,-0.0234375,-0.015625,0.0234375,-0.0078125,-0.015625,0.015625,-0.0625,0.078125,-0.0390625,-0.046875,0.015625,-0.03125,-0.03125,-0.0234375,-0.015625,0.0078125,0.0625,0.0,-0.0390625,0.0078125,-0.0078125,-0.0,0.0,-0.03125,0.0078125,0.078125,-0.03125,-0.0078125,-0.0078125,-0.0390625,0.0078125,0.0078125,-0.015625,0.0,-0.0234375,-0.0078125,0.015625,-0.0234375,-0.0234375,0.0078125,0.0,0.0078125,0.0078125,-0.0234375,-0.0,0.0,0.0078125,-0.0,0.0078125,-0.0234375,-0.015625,0.015625,-0.015625,-0.0234375,-0.015625,0.0,0.046875,0.0390625,-0.015625,-0.0234375,0.0078125,0.0234375,-0.015625,-0.0625,0.0234375,0.03125,-0.03125,-0.0078125,0.015625,0.0078125,0.015625,0.0078125,-0.015625,0.015625,0.0234375,0.0234375,-0.0078125,-0.0,-0.0,-0.0078125,-0.0,-0.0078125,0.0078125,-0.03125,-0.015625,-0.0234375,-0.0,-0.0390625,-0.03125,0.015625,-0.0,-0.0078125,-0.0078125,-0.0390625,0.0078125,0.015625,-0.015625,-0.015625,0.0,-0.0390625,0.0078125,-0.03125,-0.078125,0.0234375,0.0703125,0.0,-0.0078125,0.0234375,-0.0234375,0.015625,0.0234375,-0.0078125,0.0078125,0.0703125,0.046875,-0.0234375,-0.0078125,-0.0078125,-0.046875,0.015625,0.03125,0.0078125,-0.0546875,-0.078125,-0.03125,0.0078125,-0.0234375,0.03125,0.0234375,-0.0078125,-0.0,0.03125,0.015625,-0.0390625,-0.03125,-0.0234375,-0.046875,-0.0390625,-0.046875,-0.0234375,0.0625,0.03125,0.0,0.0,0.015625,-0.0234375,-0.0390625,-0.015625,0.0,0.046875,-0.0234375,-0.015625,0.0078125,-0.03125,-0.015625,0.0234375,0.0390625,-0.015625,-0.015625,-0.0,-0.078125,-0.0234375,-0.0078125,-0.03125,-0.03125,0.015625,0.0,0.0390625,0.03125,-0.0078125,-0.0234375,-0.0078125,-0.0234375,-0.0546875,0.015625,-0.078125,-0.03125,0.015625,0.0390625,-0.0390625,-0.0546875,-0.0234375,-0.0,-0.046875,0.0,0.0234375,-0.0234375,0.0234375,-0.0,0.015625,0.0546875,0.0234375,-0.0390625,0.0,0.046875,0.046875,0.0078125,-0.0,-0.0390625,-0.015625,-0.0390625,-0.046875,0.015625,0.0625,0.0703125,-0.0078125,-0.0078125,0.015625,0.03125,-0.0234375,-0.0234375,0.0078125,0.0390625,0.046875,-0.0234375,0.0234375,-0.0078125,-0.03125,0.0234375,0.0078125,-0.015625,0.015625,-0.0546875,-0.0390625,-0.0390625,-0.0546875,-0.046875,-0.0,-0.015625,-0.0,0.0078125,0.0,0.015625,0.0078125,0.0,-0.0078125,0.0078125,-0.0234375,-0.015625,0.0390625,0.0625,-0.0546875,0.015625,-0.0078125,0.0234375,-0.015625,0.0546875,-0.015625,0.0234375,-0.015625,-0.0,0.03125,-0.078125,0.0390625,-0.0078125,0.0390625,-0.0390625,-0.03125,0.015625,0.078125,-0.0,-0.0390625,0.015625,-0.0,-0.0078125,-0.0078125,0.0,-0.0078125,0.0078125,-0.0078125,0.0078125,-0.0,-0.0390625,-0.0625,-0.0390625,0.015625,0.0625,0.015625,0.0390625,-0.046875,0.078125,-0.078125,-0.0,0.0078125,0.078125,0.078125,-0.03125,0.0625,0.0078125,0.0234375,-0.03125,0.0390625,-0.078125,0.015625,0.03125,0.015625,0.03125,-0.0625,-0.0390625,0.0078125,-0.015625,0.0078125,0.0078125,0.0390625,-0.0,0.0390625,0.0234375,0.0625,-0.0078125,0.0,-0.03125,-0.078125,-0.0546875,-0.109375,0.046875,0.015625,0.0703125,0.0234375,0.078125,-0.0078125,-0.0234375,-0.0234375,0.0078125,-0.0234375,0.0234375,-0.0234375,-0.0234375,-0.0390625,0.03125,0.03125,0.015625,0.0078125,-0.0234375,-0.015625,0.015625,0.015625,0.03125,0.0703125,-0.03125,0.015625,0.015625,-0.0546875,-0.0234375,-0.0390625,0.0390625,-0.046875,0.0078125,-0.0078125,-0.015625,-0.0078125,-0.0625,-0.0859375,-0.03125,0.046875,-0.046875,-0.046875,0.0546875,-0.03125,0.0390625,0.0234375,-0.046875,0.0546875,0.0078125,-0.0,-0.015625,0.015625,-0.0078125,0.0,0.0078125,-0.0234375,-0.015625,-0.015625,0.0859375,0.03125,-0.015625,-0.03125,-0.03125,0.03125,0.0234375,-0.03125,-0.046875,-0.0390625,0.03125,-0.0078125,0.0,-0.015625,0.03125,0.0234375,-0.0546875,-0.0078125,-0.0234375,-0.0,-0.0546875,0.0546875,-0.0078125,0.0234375,0.0546875,-0.0625,0.015625,0.0078125,-0.0703125,-0.046875,0.0546875,0.0078125,0.015625,-0.0703125,0.03125,0.0546875,0.015625,-0.0078125,0.078125,0.0078125,-0.0703125,0.0078125,0.0,-0.0625,0.015625,-0.0,0.046875,0.078125,-0.0078125,0.03125,0.03125,-0.0390625,-0.0078125,-0.0390625,-0.1015625,0.1171875,-0.0390625,-0.0859375,0.0703125,0.046875,-0.046875,-0.015625,0.0625,0.09375,0.015625,0.0078125,-0.015625,-0.046875,-0.03125,-0.03125,0.0234375,0.03125,0.03125,0.0078125,0.0234375,-0.0234375,-0.0546875,-0.03125,0.09375,-0.015625,-0.015625,-0.0078125,0.0,0.0390625,0.0234375,-0.0078125,-0.03125,-0.03125,0.0,-0.0703125,0.0625,0.0,-0.015625,-0.0390625,-0.03125,-0.0390625,-0.0703125,0.0390625,0.0625,-0.03125,-0.0625,-0.015625,-0.046875,-0.046875,0.015625,0.015625,0.0078125,0.0,-0.0390625,-0.0078125,-0.0390625,-0.015625,-0.03125,0.0234375,0.046875,0.0,0.0078125,-0.015625,0.0703125,0.0390625,-0.0,0.0625,-0.03125,0.0078125,-0.03125,-0.046875,0.015625,0.0390625,-0.0859375,-0.0078125,-0.0546875,0.0390625,0.046875,-0.0390625,-0.0078125,-0.015625,-0.03125,0.0390625,0.0234375,0.0078125,0.0,0.03125,0.0703125,0.0,-0.015625,-0.015625,0.0,0.0,0.015625,-0.0,-0.015625,-0.0,0.0390625,-0.03125,-0.078125,-0.0234375,-0.015625,-0.0234375,-0.0390625,0.1015625,0.0859375,0.0078125,-0.0390625,0.03125,-0.015625,0.03125,-0.0234375,-0.0078125,-0.0390625,0.0234375,0.03125,-0.0078125,-0.0625,-0.078125,0.015625,0.0234375,-0.046875,-0.0390625,0.0390625,-0.0,0.0078125,0.0078125,-0.0078125,-0.0078125,0.0,0.0078125,0.0,-0.015625,0.046875,-0.0625,-0.0625,-0.03125,-0.046875,0.0625,-0.046875,-0.0625,0.0703125,-0.1015625,0.0546875,-0.0546875,-0.046875,0.015625,0.0390625,0.0390625,-0.0078125,0.0078125,-0.0390625,-0.046875,-0.0234375,0.0859375,0.0390625,-0.015625,-0.0234375,-0.015625,-0.078125,0.0078125,0.0078125,-0.015625,-0.03125,-0.015625,-0.046875,-0.046875,0.0390625,0.0390625,0.109375,-0.0,0.0625,0.0078125,-0.0703125,-0.0703125,-0.0390625,-0.015625,0.0234375,-0.0390625,0.0390625,-0.0078125,-0.0078125,-0.0390625,-0.0390625,-0.0,-0.0625,0.0078125,-0.0078125,-0.03125,-0.0078125,-0.0078125,0.0078125,0.046875,-0.0,0.0,0.0234375,-0.015625,-0.0078125,0.0234375,-0.015625,-0.1328125,0.125,-0.015625,-0.03125,-0.0078125,0.1015625,0.0234375,-0.078125,-0.015625,-0.1015625,-0.03125,0.0703125,-0.03125,-0.015625,0.0859375,0.0390625,-0.0625,0.0,-0.0390625,0.0234375,0.0,-0.0546875,0.0859375,-0.0,-0.0078125,-0.015625,0.0078125,0.0,0.015625,0.015625,0.0,0.0234375,0.0078125,0.0390625,-0.0546875,-0.0078125,0.015625,0.0234375,0.0078125,0.0078125,-0.0078125,-0.078125,0.0625,0.0703125,-0.0625,-0.078125,-0.015625,-0.0390625,0.0234375,0.0546875,-0.046875,0.046875,-0.0546875,-0.0625,-0.0703125,-0.015625,-0.0390625,0.0078125,0.1328125,-0.0234375,0.015625,-0.1328125,-0.0078125,-0.1484375,-0.0703125,0.0546875,0.0390625,0.0859375,0.0703125,0.0625,-0.0390625,0.0234375,-0.0703125,-0.0625,-0.015625,-0.0078125,0.0859375,0.03125,-0.0703125,-0.0390625,0.0625,0.0390625,0.0546875,0.0078125,0.0546875,-0.0078125,-0.0546875,-0.0390625,0.15625,-0.1015625,-0.125,0.046875,0.046875,-0.015625,0.0234375,-0.015625,0.0390625,-0.09375,-0.0078125,0.0078125,-0.1328125,0.015625,0.046875,-0.0234375,-0.0078125,0.03125,0.0234375,-0.03125,-0.078125,0.0625,0.0546875,-0.0859375,-0.0,-0.0390625,-0.0859375,-0.0625,-0.0390625,-0.03125,0.0859375,-0.015625,-0.078125,0.140625,-0.046875,-0.0,0.0546875,-0.109375,-0.1875,-0.0234375,0.015625,-0.0390625,-0.0625,0.0234375,0.1015625,-0.0,-0.0546875,0.0078125,0.03125,-0.03125,0.0859375,0.0078125,0.046875,-0.0625,0.1171875,-0.0234375,-0.109375,0.03125,-0.0625,-0.0234375,-0.0625,-0.0390625,-0.09375,0.0234375,-0.015625,0.0234375,0.0625,-0.0078125,-0.015625,0.0,0.015625,-0.0234375,0.0625,-0.0,-0.078125,0.0,-0.0859375,0.078125,0.03125,0.0390625,-0.0390625,-0.0859375,-0.03125,0.03125,0.0703125,0.0234375,-0.03125,-0.0234375,0.015625,0.0078125,0.0078125,-0.0,-0.0078125,-0.0078125,0.0078125,-0.0,-0.0078125,0.03125,-0.03125,-0.078125,-0.0546875,-0.078125,0.0078125,0.015625,-0.015625,0.03125,-0.0,-0.09375,-0.046875,0.03125,-0.03125,-0.015625,0.0234375,-0.046875,-0.0,0.0,-0.0625,0.0546875,0.140625,-0.09375,0.03125,0.0390625,0.0,-0.078125,-0.0234375,0.0,-0.0,0.0078125,0.015625,-0.015625,-0.0078125,0.0078125,-0.0,-0.0234375,-0.0390625,0.0,-0.0078125,0.0390625,-0.078125,0.015625,0.015625,0.03125,-0.0703125,0.046875,-0.046875,-0.0859375,-0.0546875,0.078125,-0.0546875,0.0078125,0.03125,0.015625,0.046875,0.0234375,0.03125,0.0078125,0.0,-0.0,-0.0703125,-0.0390625,0.046875,-0.0,-0.03125,0.0078125,0.0234375,-0.015625,-0.0234375,-0.0078125,-0.015625,0.0234375,0.046875,0.0234375,0.0234375,0.0703125,0.0078125,-0.0234375,0.0390625,0.0546875,0.0390625,-0.015625,0.0078125,0.0078125,-0.046875,-0.0234375,0.0,0.015625,0.0,-0.015625,-0.015625,-0.0234375,-0.015625,-0.0,0.0078125,-0.046875,0.015625,0.0,0.0,-0.0390625,-0.0390625,0.0703125,0.015625,0.0,-0.0390625,-0.046875,0.015625,-0.015625,-0.0390625,-0.0390625,0.046875,0.15625,-0.015625,-0.015625,-0.015625,0.0625,-0.078125,0.078125,-0.015625,-0.0859375,0.046875,-0.03125,0.0625,0.0234375,0.0234375,-0.015625,-0.0078125,-0.0078125,-0.0,0.0078125,0.0,-0.015625,0.015625,-0.0078125,-0.015625,-0.0234375,-0.0,-0.015625,-0.03125,0.0546875,-0.0,-0.0,0.0390625,-0.0390625,-0.0625,-0.0546875,0.0078125,-0.03125,0.0703125,-0.0625,-0.0234375,-0.03125,-0.0390625,-0.0078125,-0.0078125,0.0703125,0.0078125,0.0078125,0.0546875,0.09375,-0.0234375,-0.046875,-0.0859375,-0.0703125,0.0234375,0.015625,0.03125,-0.0859375,-0.0078125,0.03125,-0.0078125,-0.0625,-0.0078125,-0.0390625,-0.0,0.0078125,-0.03125,-0.0390625,-0.0390625,0.0234375,-0.03125,-0.0546875,0.015625,-0.0,-0.03125,-0.0390625,0.046875,-0.015625,0.078125,0.0234375,-0.0859375,0.046875,-0.0546875,-0.0234375,-0.0390625,-0.0234375,-0.0078125,0.015625,0.0546875,0.078125,-0.015625,0.03125,-0.0234375,-0.09375,-0.0,0.0,-0.0078125,-0.046875,-0.0078125,0.03125,-0.0703125,0.1015625,-0.0390625,-0.0859375,-0.046875,-0.015625,-0.0703125,-0.0,0.078125,0.0234375,0.03125,0.0625,0.015625,-0.03125,0.0703125,-0.0390625,-0.078125,-0.0078125,0.0234375,-0.0234375,-0.0546875,-0.09375,0.0078125,0.09375,0.0,-0.03125,-0.0234375,-0.0,-0.03125,-0.015625,-0.03125,0.03125,-0.0078125,0.0234375,-0.0546875,-0.015625,-0.078125,0.0234375,-0.015625,-0.0390625,0.015625,0.0625,-0.03125,-0.03125,-0.078125,-0.09375,-0.0390625,0.0078125,0.03125,-0.0,0.03125,-0.0078125,-0.03125,-0.046875,0.0078125,-0.015625,0.0390625,-0.03125,0.0078125,0.03125,0.0625,-0.015625,0.0625,0.015625,0.046875,0.0390625,-0.0234375,-0.0,-0.0,0.015625,0.0,-0.015625,-0.0234375,-0.0078125,0.0078125,-0.015625,-0.015625,0.0078125,-0.1171875,-0.0546875,0.046875,-0.0703125,-0.03125,-0.0703125,0.0390625,0.046875,-0.046875,-0.03125,-0.0546875,-0.0390625,-0.125,0.0703125,0.046875,0.0859375,0.1640625,-0.0546875,-0.0703125,-0.015625,0.0390625,-0.078125,0.1015625,-0.0390625,-0.0703125,-0.0703125,0.0078125,0.0,-0.0,0.0078125,0.0,-0.0078125,-0.0078125,0.0078125,-0.0,0.0234375,-0.046875,0.0625,0.15625,0.1015625,-0.078125,-0.1171875,0.015625,0.0546875,-0.0234375,-0.0703125,-0.0078125,-0.015625,-0.0546875,0.0546875,0.0078125,-0.015625,0.0,-0.0234375,-0.0390625,0.0234375,-0.046875,-0.0703125,-0.0078125,-0.046875,0.0234375,0.140625,-0.03125,-0.09375,-0.046875,-0.046875,0.03125,0.03125,0.0234375,0.0078125,0.0078125,0.046875,0.046875,0.046875,0.0390625,0.0234375,0.140625,0.03125,-0.0,0.0625,0.0234375,0.046875,0.046875,-0.015625,-0.0078125,0.0390625,0.0703125,-0.046875,-0.0390625,-0.015625,-0.0078125,0.0078125,0.0625,-0.015625,-0.03125,0.0078125,0.03125,-0.0078125,0.0390625,0.015625,-0.0,0.0546875,0.0546875,-0.0625,0.0078125,-0.03125,-0.0859375,-0.015625,-0.015625,0.0234375,-0.03125,-0.09375,-0.0078125,-0.0390625,0.0703125,0.078125,0.015625,0.03125,-0.015625,0.0546875,-0.03125,-0.09375,-0.0625,-0.0234375,-0.125,0.015625,0.0234375,-0.0,0.015625,0.0234375,0.0234375,-0.03125,0.0,-0.0078125,0.015625,0.046875,-0.0,0.0078125,-0.0625,-0.0859375,0.0234375,0.03125,0.0078125,-0.0234375,-0.0859375,-0.0234375,-0.09375,-0.109375,0.1015625,0.0625,-0.0234375,0.09375,-0.03125,-0.0390625,0.0390625,0.0390625,0.0625,-0.0078125,-0.03125,-0.0625,-0.0,0.03125,0.0234375,0.046875,-0.015625,-0.0703125,-0.0078125,-0.0390625,-0.015625,-0.0390625,-0.0234375,-0.0546875,-0.109375,0.0703125,-0.0078125,0.046875,-0.015625,-0.09375,0.0546875,-0.0390625,-0.046875,0.0546875,0.0625,-0.0390625,0.03125,-0.0078125,0.03125,-0.0078125,-0.078125,0.046875,0.1875,-0.0,-0.1796875,-0.0234375,0.0234375,-0.03125,-0.0703125,-0.0234375,0.03125,0.015625,-0.0390625,0.015625,0.0546875,0.046875,-0.03125,0.0,0.015625,-0.0390625,0.0,0.0078125,-0.046875,-0.03125,-0.0078125,-0.046875,-0.0859375,0.0078125,-0.09375,-0.0625,-0.03125,-0.0078125,0.03125,0.0078125,0.046875,-0.0078125,-0.078125,-0.1015625,0.0234375,-0.0390625,0.0390625,-0.0546875,-0.0234375,-0.078125,-0.03125,-0.1328125,-0.1015625,0.0546875,-0.0546875,-0.0859375,-0.015625,-0.015625,0.09375,0.0625,-0.0,-0.015625,-0.0390625,0.03125,-0.0390625,0.015625,0.0078125,0.046875,0.1328125,0.015625,-0.0234375,-0.0390625,0.015625,-0.1640625,0.0234375,0.0625,0.0234375,0.046875,-0.046875,-0.0078125,0.0078125,0.03125,-0.109375,-0.0390625,0.0078125,-0.0390625,-0.015625,-0.0546875,-0.1015625,-0.0390625,-0.0625,-0.0703125,-0.0703125,-0.0,-0.0078125,-0.0078125,-0.0078125,0.0078125,0.0078125,-0.0,0.0,0.0078125,-0.0078125,-0.0234375,0.015625,-0.0078125,-0.015625,0.0,-0.0,-0.0546875,0.0,-0.0078125,0.03125,-0.0234375,-0.0234375,0.0546875,-0.015625,0.015625,-0.109375,-0.0078125,-0.03125,0.0546875,-0.0546875,-0.0078125,0.1015625,-0.0234375,0.015625,0.03125,-0.046875,0.0703125,-0.0546875,-0.0625,0.0,-0.015625,0.0078125,0.015625,-0.0,0.015625,-0.015625,-0.0078125,0.015625,-0.0078125,0.03125,0.0078125,-0.0390625,0.0,-0.0859375,0.078125,-0.0,0.0546875,0.03125,-0.1328125,-0.0546875,0.03125,-0.0546875,0.0234375,-0.0,-0.0078125,0.0078125,-0.03125,-0.03125,-0.0625,0.0078125,0.125,-0.0390625,-0.0703125,0.1328125,0.0,-0.0078125,-0.046875,-0.0,-0.0234375,0.0078125,0.03125,0.03125,0.046875,0.0390625,-0.0078125,-0.015625,0.0625,-0.0234375,0.046875,-0.0625,-0.03125,0.015625,-0.015625,-0.1015625,-0.0234375,0.0234375,0.0703125,-0.078125,0.0390625,0.03125,0.0078125,0.09375,0.03125,-0.0234375,0.015625,0.046875,-0.03125,-0.015625,-0.0078125,-0.03125,-0.03125,0.09375,0.0390625,-0.0,-0.015625,-0.0078125,-0.0078125,-0.03125,-0.0078125,0.046875,0.0546875,-0.0625,0.015625,-0.015625,0.03125,0.0234375,0.0234375,-0.046875,0.046875,-0.09375,0.140625,-0.015625,-0.0546875,0.046875,0.1015625,0.0390625,-0.1015625,0.0078125,0.0078125,-0.0078125,0.0078125,0.015625,-0.0078125,0.015625,-0.0,-0.03125,-0.0078125,0.015625,-0.1015625,0.046875,-0.015625,-0.0703125,-0.0546875,-0.03125,-0.0078125,-0.0078125,-0.0078125,-0.046875,-0.0078125,0.0546875,-0.0703125,-0.015625,-0.0078125,-0.046875,-0.0390625,-0.109375,0.0078125,-0.0625,-0.03125,0.0625,0.0234375,0.0234375,-0.0703125,0.0390625,0.015625,0.015625,0.0390625,-0.0,-0.046875,0.0390625,-0.015625,-0.078125,-0.03125,0.03125,-0.015625,0.046875,-0.0,-0.0625,0.015625,-0.0859375,-0.125,0.109375,-0.015625,0.015625,-0.015625,0.03125,-0.046875,-0.0390625,0.078125,0.0703125,-0.0234375,-0.03125,0.046875,-0.078125,0.0,0.015625,-0.03125,0.0078125,0.015625,-0.0078125,-0.046875,-0.0625,0.03125,-0.0390625,0.0625,-0.0,0.015625,0.015625,0.046875,-0.0078125,-0.046875,0.0,0.015625,0.0,-0.03125,-0.0390625,0.0546875,0.046875,0.03125,0.0546875,0.0546875,0.0234375,-0.0625,-0.0390625,0.0546875,0.03125,0.046875,0.0703125,-0.0546875,0.0,-0.03125,0.0078125,-0.0625,-0.03125,0.0546875,0.015625,-0.0,0.03125,0.0078125,0.0078125,-0.0390625,-0.0859375,-0.0625,0.015625,0.015625,0.0390625,0.0546875,0.03125,-0.0078125,-0.078125,0.046875,-0.09375,0.0546875,0.0078125,0.0546875,0.0625,0.0234375,-0.015625,-0.015625,0.0078125,-0.03125,-0.0703125,-0.015625,-0.046875,-0.109375,0.015625,0.015625,0.0,-0.0390625,0.03125,0.0625,0.0859375,-0.0234375,0.03125,-0.0234375,0.0078125,0.046875,-0.0625,-0.03125,0.046875,0.0078125,-0.015625,-0.015625,0.0,-0.0,0.0078125,-0.0078125,0.0078125,-0.0,0.03125,0.015625,0.015625,-0.046875,-0.0703125,-0.015625,-0.015625,-0.0078125,-0.0,0.0859375,0.0078125,0.0078125,0.0625,0.0390625,-0.046875,0.0078125,0.0078125,0.015625,0.0078125,-0.046875,-0.0546875,-0.0078125,-0.0546875,-0.03125,-0.0625,-0.109375,0.125,0.1015625,-0.0078125,0.0,0.0078125,0.0078125,-0.0078125,-0.015625,0.0,-0.015625,0.0078125,-0.1015625,-0.0234375,0.0625,-0.015625,-0.046875,0.1171875,0.0546875,-0.09375,0.0546875,0.03125,-0.046875,0.046875,-0.0078125,0.09375,-0.1015625,0.0078125,-0.0,0.0078125,-0.0,0.0625,-0.03125,-0.0859375,0.0859375,-0.09375,-0.0859375,0.0859375,-0.0625,0.0546875,0.046875,-0.0234375,-0.0234375,-0.0078125,-0.03125,0.0234375,0.046875,0.0078125,-0.0234375,-0.0078125,-0.0390625,-0.0234375,-0.03125,-0.03125,0.015625,-0.0234375,0.046875,-0.0234375,-0.0390625,-0.03125,0.015625,0.0,-0.03125,0.0390625,0.0,0.0234375,-0.0078125,-0.015625,-0.0078125,0.0078125,0.0,-0.0234375,0.03125,0.015625,0.0078125,0.0078125,-0.0234375,0.015625,-0.0546875,0.015625,0.0234375,-0.046875,-0.0234375,0.03125,-0.015625,0.0078125,-0.0078125,-0.0078125,-0.1015625,-0.0546875,0.0390625,0.015625,0.0546875,-0.0234375,-0.0625,-0.03125,0.03125,-0.015625,0.0625,-0.0625,-0.046875,0.09375,-0.0078125,0.0,-0.015625,0.0,0.0078125,0.0,-0.0078125,0.0078125,0.0390625,0.0234375,0.0078125,-0.0546875,0.03125,0.015625,-0.0625,0.0625,-0.015625,0.0234375,0.0703125,-0.0390625,0.0234375,-0.0234375,0.0078125,-0.0546875,-0.0234375,-0.09375,0.0546875,0.0078125,0.0390625,0.0078125,0.0078125,-0.0,-0.0234375,-0.015625,-0.0625,0.0546875,0.0859375,-0.0546875,-0.015625,-0.015625,-0.0859375,-0.078125,0.1015625,-0.0078125,0.0859375,0.0625,0.0234375,-0.078125,0.0390625,-0.078125,-0.0625,-0.0078125,0.046875,-0.015625,-0.0234375,-0.0546875,-0.03125,-0.046875,0.0078125,-0.015625,-0.0,-0.0625,0.1015625,0.0625,-0.0703125,0.0703125,-0.015625,-0.0390625,0.0078125,0.0,-0.0703125,0.0,-0.0078125,0.015625,-0.0703125,-0.0390625,0.0546875,-0.0390625,0.015625,0.0234375,0.0390625,-0.0234375,-0.03125,0.03125,-0.0625,-0.0234375,-0.0078125,-0.015625,-0.015625,0.0859375,0.03125,-0.0546875,-0.046875,0.0234375,-0.0703125,-0.0703125,0.046875,0.0078125,0.03125,-0.0078125,-0.015625,-0.046875,-0.109375,-0.0625,0.109375,-0.015625,0.0078125,-0.046875,0.0625,-0.0234375,0.0078125,-0.046875,-0.0,-0.0390625,0.0078125,0.0234375,-0.03125,0.0078125,-0.046875,0.0078125,-0.078125,0.0078125,0.03125,0.0625,-0.0625,0.046875,0.0390625,-0.078125,0.0625,0.015625,0.0234375,-0.0546875,-0.0078125,-0.0078125,0.03125,0.046875,-0.03125,-0.0078125,-0.0546875,0.015625,0.0546875,0.015625,-0.015625,0.0234375,-0.0234375,0.078125,0.03125,-0.0234375,-0.09375,0.0078125,-0.015625,-0.0078125,-0.015625,-0.0078125,-0.015625,-0.0078125,-0.015625,-0.0234375,0.0234375,-0.0,-0.0078125,-0.0,0.0078125,0.0703125,0.0078125,0.0078125,-0.0703125,-0.0390625,0.03125,-0.046875,-0.0,0.0078125,-0.0234375,0.0078125,0.0234375,-0.046875,-0.1015625,0.046875,0.0078125,0.0234375,0.0234375,0.0,0.0234375,0.0234375,0.03125,0.015625,-0.0390625,0.0078125,-0.015625,0.0078125,-0.015625,-0.0,0.015625,-0.0078125,-0.0078125,0.0,-0.0,0.0078125,-0.0234375,0.0078125,0.0390625,-0.03125,-0.0234375,-0.03125,0.0078125,-0.0078125,-0.0390625,-0.046875,-0.0859375,0.0078125,0.0546875,0.0078125,-0.0390625,-0.0078125,0.0,0.0625,-0.03125,0.03125,0.0,0.046875,0.0,0.015625,-0.046875,-0.0546875,-0.0390625,0.0546875,-0.0234375,-0.0,0.015625,-0.0234375,-0.03125,-0.015625,-0.015625,-0.015625,-0.0625,-0.0078125,0.0703125,-0.0390625,-0.0625,-0.0625,-0.046875,0.0078125,-0.03125,-0.015625,0.015625,0.0546875,0.0078125,-0.0546875,0.03125,-0.0078125,-0.0078125,0.0390625,-0.03125,-0.046875,-0.015625,-0.0078125,0.03125,0.015625,0.0,0.0390625,0.0546875,-0.0078125,0.0078125,-0.0546875,-0.015625,0.09375,-0.03125,-0.0078125,0.0,-0.03125,0.0546875,0.0234375,0.0,0.0625,-0.015625,-0.0078125,-0.03125,-0.0390625,-0.03125,0.015625,-0.0390625,-0.0234375,-0.015625,0.0625,0.0,-0.015625,0.0078125,0.0078125,-0.015625,0.0,0.0234375,0.0234375,0.0234375,0.03125,-0.0078125,-0.0,0.0078125,-0.015625,-0.0,0.015625,-0.0390625,0.0078125,-0.0390625,0.0390625,0.015625,-0.03125,-0.015625,0.0390625,0.1484375,0.0234375,-0.0859375,0.015625,-0.015625,-0.0,-0.046875,-0.015625,0.03125,0.0078125,0.015625,-0.0390625,0.0390625,-0.0390625,-0.046875,-0.046875,-0.0390625,-0.0390625,0.1484375,0.015625,0.0546875,0.0625,-0.0390625,-0.0234375,0.0234375,0.1015625,0.03125,-0.0078125,-0.0390625,-0.0234375,0.0546875,-0.015625,0.0234375,0.015625,0.0390625,0.015625,0.0,-0.046875,0.0078125,0.0078125,0.0078125,-0.0546875,0.0078125,-0.046875,-0.0859375,0.0234375,-0.015625,0.0234375,0.046875,-0.0234375,-0.0859375,-0.0625,-0.015625,-0.015625,0.0078125,-0.046875,0.03125,0.0390625,-0.015625,-0.0703125,-0.046875,0.0234375,-0.0078125,0.0234375,0.0078125,-0.0234375,0.03125,-0.0078125,0.0234375,0.0625,-0.015625,0.0546875,0.0234375,-0.0390625,-0.0234375,-0.046875,-0.03125,0.0625,0.046875,0.0234375,-0.1171875,0.0859375,-0.046875,0.0703125,-0.015625,0.015625,0.0078125,0.0234375,-0.015625,0.0,0.1640625,0.03125,-0.0859375,-0.0859375,0.0,0.03125,-0.015625,0.0078125,0.0078125,0.0625,-0.0546875,-0.0078125,-0.109375,0.078125,0.015625,0.0078125,-0.03125,-0.015625,0.0,-0.0234375,-0.015625,-0.046875,-0.0078125,0.015625,0.015625,-0.03125,-0.0859375,0.015625,-0.0078125,0.0,0.015625,-0.0078125,0.0,0.0234375,-0.0234375,0.015625,-0.0078125,0.0234375,-0.0078125,0.0,-0.0234375,0.046875,-0.03125,0.0078125,0.0,-0.0078125,-0.0078125,0.0,0.0078125,0.015625,0.0,0.0,-0.0078125,-0.0390625,0.0,-0.0859375,0.0546875,-0.015625,0.0859375,-0.0234375,-0.015625,-0.0,-0.0078125,0.0078125,-0.0234375,0.0390625,-0.0078125,0.03125,-0.0703125,-0.0625,0.0,-0.0078125,-0.0078125,-0.078125,-0.0078125,-0.03125,0.0859375,0.015625,-0.0,-0.0,0.0,-0.0,0.0078125,-0.0078125,-0.0,0.0,-0.015625,0.0,-0.015625,-0.0,0.0,-0.1015625,0.015625,-0.0234375,-0.03125,-0.015625,-0.015625,0.046875,0.0078125,-0.0234375,0.1875,-0.1015625,-0.0078125,0.0546875,-0.0078125,-0.0390625,0.0390625,0.0546875,-0.015625,0.0078125,-0.0,-0.03125,-0.0703125,-0.0234375,-0.0703125,-0.046875,0.0078125,0.0078125,0.015625,-0.0703125,-0.03125,0.0,-0.046875,-0.0,0.0,0.0234375,-0.0078125,0.0,-0.0625,-0.0,-0.0390625,-0.0625,0.0078125,-0.03125,0.0,0.0,0.078125,-0.015625,-0.0078125,-0.015625,-0.0078125,0.0078125,0.015625,-0.0078125,0.0,0.03125,-0.0078125,-0.0,-0.0078125,-0.03125,-0.015625,-0.0078125,-0.0078125,0.0078125,-0.0,-0.0390625,-0.0078125,0.015625,-0.0,-0.015625,-0.0234375,-0.0390625,-0.0,-0.09375,-0.140625,0.0,0.015625,0.03125,-0.0078125,0.0078125,0.0546875,-0.015625,-0.0078125,0.0078125,-0.046875,-0.1640625,0.046875,-0.0234375,-0.0078125,0.0078125,-0.0078125,0.0,0.015625,0.0,0.0078125,0.0078125,-0.015625,-0.015625,-0.0078125,0.015625,-0.015625,-0.03125,0.0234375,-0.015625,0.0390625,0.0,-0.0234375,-0.0234375,0.0,-0.0390625,0.03125,-0.015625,0.0859375,-0.09375,-0.046875,-0.0,-0.0078125,0.015625,-0.015625,-0.09375,-0.0390625,0.1484375,-0.09375,0.0078125,-0.015625,-0.046875,0.0078125,-0.0234375,-0.046875,-0.0390625,0.0,0.03125,-0.0234375,-0.0625,-0.0234375,0.015625,-0.0546875,-0.0625,-0.015625,-0.0546875,0.03125,-0.03125,0.0078125,-0.0234375,-0.015625,-0.0625,0.0703125,-0.03125,0.015625,-0.0703125,-0.0,0.0078125,-0.03125,0.0234375,-0.03125,-0.0390625,-0.015625,0.1015625,-0.0546875,-0.0390625,-0.046875,-0.0078125,-0.0078125,0.046875,-0.0078125,-0.015625,0.0390625,0.0390625,-0.015625,-0.0078125,0.0,0.0234375,-0.015625,-0.0390625,0.0,-0.0,0.015625,-0.015625,-0.0078125,-0.0234375,0.0078125,0.15625,0.0078125,-0.0,-0.03125,-0.0859375,-0.03125,-0.0078125,-0.0234375,-0.0078125,-0.046875,0.0703125,-0.0703125,-0.0,0.03125,-0.0078125,-0.046875,-0.0703125,0.0,-0.0234375,0.0078125,-0.046875,-0.0234375,-0.03125,-0.0234375,-0.0078125,-0.03125,-0.0078125,0.03125,0.0625,-0.0,-0.015625,-0.0078125,-0.015625,0.0625,-0.015625,-0.03125,0.0546875,-0.09375,-0.03125,0.0390625,-0.0078125,-0.015625,-0.0078125,-0.0078125,0.0078125,-0.078125,0.0703125,-0.0,0.0625,-0.015625,-0.0234375,0.03125,0.0,0.0625,-0.0078125,-0.0078125,-0.0234375,-0.0390625,-0.1015625,-0.046875,-0.0078125,-0.015625,0.0078125,0.0078125,0.015625,-0.0,-0.0078125,0.0234375,-0.0078125,0.0,-0.0078125,0.0078125,0.1015625,-0.046875,0.0546875,0.0625,-0.0859375,-0.09375,-0.0546875,-0.0234375,-0.0234375,-0.0234375,0.0,0.0390625,0.046875,0.03125,0.046875,-0.0078125,-0.0078125,-0.0390625,-0.0390625,0.0078125,-0.03125,-0.03125,-0.0,0.1015625,0.0,0.015625,0.0,-0.0078125,-0.0078125,-0.0078125,-0.0078125,-0.0078125,0.0078125,-0.015625,0.0234375,-0.0703125,-0.0078125,-0.1171875,0.0703125,0.1015625,0.0390625,-0.078125,0.0859375,-0.03125,0.140625,-0.015625,-0.0625,-0.0859375,0.0703125,0.015625,-0.0,0.0546875,0.03125,-0.0078125,0.0,0.015625,0.015625,-0.0078125,-0.078125,0.0234375,0.03125,-0.03125,-0.046875,0.0546875,0.0546875,-0.03125,0.0234375,-0.0703125,-0.03125,-0.015625,-0.0546875,-0.0078125,-0.0234375,-0.046875,-0.046875,-0.015625,0.109375,0.0546875,-0.0078125,-0.0546875,0.0,-0.0,-0.015625,0.0390625,-0.0078125,0.0078125,0.0078125,0.0546875,0.03125,0.015625,-0.0390625,-0.0078125,-0.0078125,-0.0,-0.0390625,-0.015625,-0.0078125,0.0078125,-0.0078125,-0.0390625,0.0078125,-0.015625,0.0859375,0.0703125,-0.03125,0.015625,-0.015625,-0.03125,-0.0546875,0.0625,-0.0703125,0.0078125,0.015625,-0.0546875,0.0078125,-0.0234375,-0.0234375,-0.0078125,0.0,0.03125,0.0078125,-0.0625,-0.0703125,0.015625,0.0078125,-0.0078125,-0.0078125,0.0078125,-0.015625,-0.0,0.0,0.0234375,-0.03125,0.03125,0.03125,0.046875,-0.03125,-0.0078125,-0.0234375,0.0078125,-0.0078125,0.0078125,0.0,0.015625,-0.0390625,-0.0859375,0.046875,0.0234375,0.0234375,-0.0390625,0.0390625,-0.0,-0.046875,0.0390625,-0.078125,0.015625,0.03125,-0.0390625,-0.0234375,0.0078125,-0.0078125,-0.03125,0.03125,0.1171875,0.0234375,-0.0625,0.0078125,-0.015625,0.0390625,-0.046875,-0.0078125,0.0234375,-0.03125,-0.015625,-0.0,-0.015625,0.03125,0.0,-0.0546875,-0.0,0.0234375,-0.0078125,0.078125,-0.046875,-0.078125,0.0078125,0.0078125,-0.046875,-0.03125,-0.140625,-0.0,0.1015625,0.015625,-0.0859375,0.09375,-0.015625,-0.046875,-0.0234375,0.046875,-0.0078125,-0.0546875,0.0078125,-0.0390625,-0.0078125,0.03125,-0.015625,0.0390625,-0.0,-0.0078125,-0.03125,-0.0078125,-0.0078125,-0.015625,0.09375,0.0703125,0.1015625,-0.03125,-0.03125,-0.0,0.0546875,-0.015625,0.046875,0.015625,0.015625,-0.0390625,-0.0625,-0.0234375,-0.0546875,0.09375,0.0078125,-0.0,-0.0390625,-0.0625,-0.0390625,-0.03125,-0.09375,-0.0078125,-0.0546875,0.078125,0.0234375,-0.0078125,0.015625,-0.0390625,0.03125,-0.0859375,0.0234375,0.078125,0.0390625,-0.0546875,-0.0078125,0.03125,-0.0390625,0.046875,-0.015625,0.0390625,-0.0703125,0.0390625,0.03125,0.0078125,0.078125,0.0703125,-0.0625,-0.0546875,-0.0390625,-0.046875,-0.1171875,0.0234375,-0.0703125,-0.015625,-0.0234375,-0.015625,0.03125,-0.0078125,0.0234375,0.0234375,0.0,-0.015625,-0.0078125,-0.015625,-0.015625,0.0078125,0.0078125,-0.0,-0.0,0.0078125,0.0390625,-0.0859375,0.0390625,0.0078125,-0.078125,0.0078125,0.0234375,-0.03125,0.0859375,0.0,-0.03125,0.0078125,0.0859375,-0.09375,-0.046875,0.078125,-0.078125,0.109375,-0.0703125,-0.046875,-0.0546875,-0.0625,-0.0234375,0.015625,-0.1171875,0.15625,-0.0,0.0078125,0.0078125,-0.0078125,0.0078125,0.0078125,-0.0078125,-0.0,0.0078125,0.0,-0.0390625,-0.0546875,-0.0,-0.0078125,-0.1328125,0.1328125,0.0546875,-0.078125,0.078125,0.0625,-0.1015625,0.1171875,0.0390625,-0.1171875,-0.0078125,-0.0625,0.0625,-0.0,-0.0234375,0.0859375,0.09375,-0.0390625,0.1640625,-0.109375,0.0390625,0.0703125,-0.0390625,0.0078125,-0.0078125,0.03125,0.0234375,-0.0234375,-0.0234375,-0.0703125,-0.0078125,-0.03125,0.0078125,0.0546875,-0.015625,0.0078125,0.0078125,-0.0,-0.0,-0.0234375,0.0078125,0.0078125,-0.078125,-0.0078125,-0.015625,-0.046875,0.0078125,0.015625,0.0078125,0.0,-0.03125,-0.0390625,-0.0078125,0.015625,-0.0625,0.0234375,0.03125,0.015625,-0.0,-0.0234375,-0.0390625,0.0078125,-0.0703125,0.078125,-0.0625,0.03125,0.0390625,-0.0,-0.0234375,0.046875,-0.0390625,-0.0625,-0.0390625,-0.0234375,0.0625,0.0,0.015625,-0.046875,0.03125,-0.046875,0.0234375,-0.03125,0.0546875,-0.09375,0.046875,-0.0390625,0.0078125,0.0078125,-0.015625,-0.015625,0.0,-0.03125,-0.015625,0.015625,0.0234375,0.0390625,-0.0234375,0.046875,0.0234375,0.03125,-0.0078125,0.0546875,-0.0,0.0625,0.09375,-0.0390625,0.0625,-0.0078125,-0.0234375,-0.0859375,0.0078125,-0.0390625,-0.0234375,0.0234375,-0.015625,0.0234375,-0.03125,0.03125,-0.0625,-0.015625,0.03125,-0.0390625,0.0,-0.0703125,0.015625,-0.015625,-0.0390625,-0.0546875,-0.0546875,0.0234375,0.0234375,-0.015625,-0.0859375,0.0078125,-0.0703125,-0.0703125,0.046875,-0.15625,0.1875,-0.09375,0.0234375,-0.0234375,-0.0078125,0.0625,0.046875,-0.0390625,0.0859375,-0.078125,0.03125,0.0625,0.015625,0.03125,-0.0,-0.0078125,-0.078125,-0.0390625,-0.0625,0.0234375,-0.0703125,0.046875,0.0390625,-0.0703125,0.0546875,0.0390625,0.078125,0.0078125,0.109375,0.015625,0.078125,0.0234375,0.015625,-0.0703125,-0.015625,-0.03125,0.078125,-0.0078125,0.0234375,-0.0234375,-0.0,0.0,0.046875,0.015625,-0.0703125,0.140625,-0.0,0.015625,0.0703125,0.046875,-0.015625,0.0390625,-0.0234375,-0.0234375,-0.0625,-0.0234375,-0.0390625,-0.03125,-0.0859375,-0.0703125,-0.046875,-0.0234375,-0.09375,0.03125,-0.0,0.015625,-0.0546875,-0.0078125,-0.046875,-0.140625,-0.1171875,-0.0078125,0.015625,-0.0234375,-0.03125,-0.140625,-0.015625,0.015625,-0.0390625,-0.0546875,-0.015625,-0.046875,0.0703125,0.0859375,0.0234375,0.0078125,-0.0625,-0.0390625,0.0390625,0.03125,0.0546875,-0.0234375,0.0078125,0.203125,-0.0,-0.1015625,0.03125,-0.0390625,-0.0546875,-0.0546875,0.0,0.015625,-0.0078125,0.0078125,0.0078125,0.015625,-0.0234375,-0.0078125,0.0078125,-0.0,0.0546875,0.0390625,-0.0078125,-0.078125,-0.1015625,-0.0546875,-0.0,-0.0703125,0.03125,-0.046875,-0.015625,0.0703125,0.0625,-0.046875,0.0078125,0.0078125,-0.0390625,-0.0,-0.046875,-0.0625,-0.0625,-0.03125,0.046875,-0.046875,-0.0078125,0.0078125,-0.0078125,0.015625,-0.0078125,0.0078125,-0.0078125,0.0078125,0.0078125,0.0078125,-0.0078125,-0.0,-0.0703125,-0.0390625,0.0234375,-0.0546875,0.0234375,-0.0234375,-0.0703125,0.0,-0.0703125,-0.03125,-0.0390625,-0.046875,-0.09375,0.015625,0.046875,0.0546875,0.046875,0.0078125,0.09375,-0.0078125,0.03125,0.03125,-0.0859375,0.015625,-0.046875,-0.0625,0.0078125,-0.0078125,-0.078125,-0.0078125,-0.046875,0.03125,0.0078125,-0.0390625,0.0234375,0.015625,-0.015625,0.0859375,-0.0078125,-0.0078125,0.0078125,0.1171875,0.015625,-0.0390625,0.0078125,-0.0,-0.015625,-0.0078125,-0.0234375,-0.015625,-0.0625,-0.046875,-0.015625,-0.0546875,0.0234375,-0.0234375,0.0234375,-0.0234375,-0.0546875,0.0078125,0.015625,0.0078125,0.0078125,-0.0234375,-0.03125,0.015625,0.0078125,-0.046875,-0.0390625,0.0078125,0.03125,-0.0546875,0.015625,-0.046875,0.03125,-0.1171875,0.046875,-0.0625,-0.015625,0.015625,0.03125,0.0703125,0.0078125,-0.046875,0.09375,-0.046875,0.03125,-0.03125,-0.015625,0.0859375,-0.0078125,-0.0234375,-0.0,0.03125,0.0390625,0.0,0.03125,0.015625,0.0078125,-0.015625,-0.015625,-0.0234375,-0.0625,-0.0078125,-0.03125,-0.015625,-0.0078125,0.0234375,0.0546875,0.0546875,0.03125,0.0234375,-0.03125,-0.078125,0.0390625,0.078125,0.03125,-0.0078125,0.015625,-0.0,-0.109375,0.046875,-0.078125,-0.0859375,-0.0546875,-0.046875,0.0546875,0.0234375,0.0703125,-0.09375,0.109375,-0.1171875,0.03125,-0.0390625,-0.0078125,0.015625,-0.0546875,0.0234375,0.0390625,-0.0078125,0.0703125,0.0546875,-0.078125,0.0546875,0.03125,0.0078125,0.0703125,-0.0,-0.03125,0.015625,-0.0078125,-0.046875,0.015625,0.09375,-0.0390625,0.0390625,-0.0390625,-0.1171875,-0.0859375,0.0078125,0.0859375,0.0546875,0.0390625,0.0390625,-0.0078125,-0.0078125,0.0703125,-0.0625,0.0,-0.046875,0.0234375,0.0625,-0.0234375,0.046875,0.015625,0.015625,-0.0546875,0.0234375,0.046875,0.0078125,-0.0078125,-0.0234375,-0.0078125,0.0078125,-0.015625,-0.015625,-0.0234375,0.0078125,-0.03125,0.015625,-0.046875,0.0625,-0.03125,-0.015625,0.046875,-0.0546875,-0.1328125,-0.0078125,0.0,-0.1171875,-0.0546875,-0.015625,0.0,-0.0546875,0.0625,0.1796875,0.0078125,-0.0,0.0,0.03125,0.0,-0.0546875,0.09375,-0.0703125,0.0390625,-0.0390625,0.03125,0.015625,0.046875,-0.0703125,-0.0,-0.046875,0.046875,0.0390625,0.0703125,0.078125,-0.03125,0.046875,-0.0,-0.0703125,0.0390625,-0.1015625,-0.0625,-0.0234375,0.0546875,-0.0234375,-0.0390625,0.0234375,0.015625,0.0234375,-0.015625,-0.0,-0.015625,-0.015625,0.0078125,-0.015625,0.0,-0.0,-0.0078125,-0.015625,-0.0,-0.0,-0.0234375,-0.015625,0.015625,-0.0546875,-0.0390625,-0.0703125,0.109375,-0.03125,-0.0546875,-0.03125,-0.0546875,-0.03125,0.0234375,-0.0390625,-0.015625,0.015625,0.03125,-0.015625,0.015625,-0.03125,-0.03125,0.0546875,-0.0,0.0625,0.046875,-0.0625,-0.015625,0.0,-0.0,0.0078125,-0.0,-0.0078125,0.015625,-0.0078125,-0.0,-0.0078125,-0.0546875,-0.046875,-0.0546875,-0.015625,-0.1015625,0.0625,0.0625,-0.0859375,0.078125,-0.0546875,-0.015625,0.0078125,-0.0,0.0390625,-0.0078125,-0.0703125,0.015625,0.015625,0.0234375,-0.046875,-0.0078125,0.1328125,0.0625,0.0703125,0.015625,-0.125,-0.0625,0.0234375,-0.0,0.015625,0.015625,0.0390625,-0.0234375,0.0703125,0.0546875,-0.03125,0.0078125,0.0234375,0.015625,0.03125,-0.0234375,-0.0390625,-0.0234375,-0.0390625,0.0546875,0.015625,-0.0234375,-0.0234375,-0.0234375,-0.0625,-0.046875,-0.0234375,-0.0390625,0.0078125,-0.0078125,-0.015625,-0.03125,0.015625,0.0,-0.0078125,0.0078125,0.015625,-0.0,0.0,-0.0234375,-0.0,-0.015625,0.0078125,0.0078125,-0.046875,-0.0625,-0.03125,0.0390625,0.1015625,-0.0546875,0.0,-0.0546875,-0.0703125,-0.0546875,0.0390625,0.0234375,0.0078125,0.0,-0.046875,-0.0234375,-0.0,0.0625,-0.0078125,-0.0078125,0.0390625,-0.0,0.0,-0.0234375,-0.0,-0.015625,0.0,-0.015625,-0.015625,-0.0078125,0.0546875,0.0,0.0234375,0.0078125,0.046875,-0.0546875,0.0078125,0.0078125,-0.0078125,-0.0234375,0.0546875,-0.1015625,0.03125,-0.015625,-0.03125,-0.015625,0.0390625,-0.03125,-0.0625,-0.015625,-0.015625,-0.0234375,0.0390625,-0.0078125,-0.03125,0.109375,0.0546875,-0.0234375,0.0390625,-0.03125,-0.0390625,-0.1015625,0.0078125,0.0078125,-0.015625,0.0078125,-0.0546875,-0.015625,-0.03125,0.015625,0.0390625,-0.03125,0.0703125,-0.0234375,0.0546875,-0.015625,0.109375,-0.046875,-0.0703125,-0.0625,0.0,0.0078125,0.0,-0.0546875,0.0390625,-0.015625,-0.0625,-0.1015625,0.078125,-0.0234375,-0.0546875,0.015625,-0.046875,0.0859375,0.0078125,0.046875,0.015625,0.03125,0.0234375,0.0234375,-0.0546875,-0.0078125,-0.015625,0.015625,0.0390625,-0.0546875,-0.046875,0.0078125,-0.015625,0.0390625,0.0390625,0.015625,-0.046875,-0.0234375,0.0078125,-0.0234375,-0.015625,0.015625,-0.0078125,-0.0078125,0.0,-0.03125,0.0390625,-0.015625,0.0,-0.0546875,-0.0546875,-0.046875,0.0078125,-0.09375,0.0390625,-0.0078125,0.015625,0.0234375,0.0546875,0.046875,-0.03125,0.0234375,-0.0703125,0.1171875,0.0078125,-0.046875,-0.078125,-0.015625,-0.03125,-0.015625,0.0390625,-0.015625,0.0234375,-0.03125,-0.03125,-0.0234375,0.0390625,0.015625,0.015625,-0.0234375,-0.03125,0.03125,-0.0625,-0.0546875,0.0234375,-0.0546875,0.03125,-0.0546875,0.0078125,0.0390625,0.125,-0.015625,0.0078125,-0.0078125,0.03125,-0.0859375,-0.0390625,-0.0078125,0.015625,-0.0078125,0.0,-0.015625,0.0078125,0.0078125,-0.0078125,0.015625,-0.0,0.078125,0.0859375,0.0,-0.0859375,-0.0703125,-0.0390625,-0.0234375,-0.03125,0.0078125,0.0234375,0.0234375,0.0703125,-0.0625,0.015625,-0.0859375,0.0625,0.015625,0.0546875,-0.0078125,-0.0234375,0.046875,0.0,-0.0390625,-0.015625,-0.015625,-0.0234375,0.0078125,-0.0078125,0.0234375,0.0078125,-0.0,-0.0078125,0.0,0.0,0.015625,0.0078125,0.0703125,-0.0625,0.078125,0.0,-0.0234375,0.109375,0.03125,-0.0078125,0.0390625,-0.03125,-0.0546875,-0.03125,-0.0390625,0.03125,-0.0625,0.0078125,0.0078125,0.0390625,-0.0078125,-0.015625,-0.0078125,-0.015625,0.0546875,-0.0625,0.0625,0.109375,0.0390625,0.0234375,0.0390625,0.0,-0.0546875,-0.0546875,0.0625,0.0234375,0.0078125,0.0234375,-0.03125,-0.015625,-0.0546875,-0.015625,0.0,-0.046875,-0.0234375,-0.1484375,-0.0078125,0.0078125,-0.0234375,-0.0546875,0.0,0.015625,-0.0078125,-0.0078125,0.015625,-0.0390625,-0.015625,-0.0546875,-0.0390625,0.015625,0.0546875,0.0078125,-0.0,0.0078125,0.0390625,-0.0234375,0.0078125,-0.03125,-0.0625,0.0078125,-0.0390625,-0.03125,0.015625,-0.0078125,-0.046875,0.0234375,-0.0625,0.0625,-0.078125,-0.0234375,0.0078125,-0.0390625,0.015625,-0.0546875,-0.0234375,-0.03125,0.046875,0.0,0.0703125,-0.0078125,0.03125,-0.03125,0.0,0.0,0.0078125,-0.0,-0.0078125,0.0,0.0234375,0.03125,0.0234375,0.015625,-0.015625,-0.0703125,-0.0625,-0.0625,0.015625,0.0390625,-0.0078125,0.0078125,0.046875,-0.0,0.046875,0.03125,-0.015625,0.046875,-0.0234375,-0.0390625,0.015625,0.0,0.015625,0.0,0.03125,-0.0546875,0.015625,0.0546875,-0.0546875,0.015625,-0.0625,0.046875,-0.015625,-0.09375,0.0078125,-0.1015625,0.03125,-0.015625,0.046875,-0.0,-0.0390625,-0.1171875,0.0390625,-0.078125,0.0234375,0.0234375,0.0,0.015625,0.03125,0.0859375,0.0546875,-0.0859375,-0.0625,-0.0234375,0.0078125,-0.0625,0.0546875,0.015625,-0.046875,0.0390625,-0.03125,0.03125,-0.0234375,-0.0078125,0.046875,-0.0078125,-0.0,0.0078125,-0.0078125,-0.0234375,-0.03125,0.015625,-0.0234375,0.046875,0.0390625,-0.078125,-0.0078125,-0.03125,-0.0078125,0.015625,-0.0859375,0.0234375,0.0859375,0.0,0.03125,-0.0390625,0.0,0.03125,-0.0390625,-0.015625,0.03125,0.09375,0.03125,-0.0703125,-0.0625,-0.0078125,0.0546875,0.0546875,0.015625,-0.0,0.109375,-0.0390625,-0.078125,0.0703125,-0.046875,0.0625,0.0234375,-0.0703125,-0.03125,-0.0859375,0.0078125,0.0,-0.0,0.03125,-0.015625,-0.140625,-0.0625,0.09375,-0.140625,0.1328125,-0.0234375,0.0234375,-0.0078125,-0.0703125,-0.0078125,0.0234375,-0.0234375,0.015625,0.078125,-0.0078125,0.03125,0.0078125,0.0703125,-0.078125,0.0390625,0.0078125,-0.0,-0.078125,0.0390625,0.125,0.0546875,-0.0234375,-0.0390625,0.0,0.046875,-0.03125,-0.0390625,0.0078125,0.0078125,-0.0078125,-0.0078125,0.0078125,-0.015625,-0.0078125,-0.0078125,-0.015625,-0.0703125,-0.015625,0.03125,0.0703125,-0.0390625,-0.015625,-0.015625,0.0078125,-0.0234375,-0.015625,0.0078125,-0.0234375,-0.015625,0.015625,-0.0078125,0.0078125,0.0078125,-0.03125,-0.0078125,0.015625,-0.0234375,-0.0390625,-0.0625,-0.03125,0.0234375,0.015625,-0.0390625,-0.0078125,0.0234375,-0.0,-0.0078125,0.0078125,0.015625,-0.0078125,-0.0078125,-0.0078125,0.03125,0.046875,-0.03125,-0.0234375,0.0390625,-0.0625,0.046875,-0.0,-0.0390625,0.0,0.078125,-0.0546875,-0.015625,-0.0546875,-0.0703125,0.015625,0.0234375,-0.0234375,0.015625,0.0234375,-0.0078125,-0.046875,-0.0078125,-0.03125,0.0390625,0.0703125,-0.015625,-0.0078125,-0.0,0.0546875,0.0234375,-0.015625,0.03125,-0.0,0.0,-0.0078125,0.0078125,-0.0234375,0.0234375,0.0078125,-0.0625,-0.0390625,0.0703125,-0.0078125,-0.03125,-0.015625,0.0078125,-0.0078125,-0.0234375,-0.0234375,-0.0234375,-0.015625,-0.015625,-0.03125,-0.0078125,0.0078125,-0.015625,-0.015625,-0.015625,-0.0078125,0.0234375,0.0,-0.0078125,-0.0078125,0.0,-0.0078125,-0.0234375,0.015625,-0.0,0.0234375,0.0,0.03125,-0.0625,-0.0703125,0.0546875,0.0859375,-0.0234375,0.0859375,0.078125,0.0234375,-0.0078125,0.03125,0.015625,-0.0625,-0.0625,0.0390625,-0.0078125,0.046875,0.0390625,-0.0390625,0.0,-0.0,0.0,0.0,0.0078125,0.0,-0.03125,0.0234375,0.0234375,0.015625,0.015625,0.0078125,-0.015625,-0.0078125,-0.0234375,0.0,-0.0234375,-0.0078125,-0.0234375,-0.0546875,-0.0390625,0.0,-0.015625,0.03125,0.015625,0.0,-0.0,0.0078125,0.0234375,0.109375,0.0546875,-0.046875,-0.0,0.03125,-0.0546875,-0.03125,-0.0625,-0.0625,-0.015625,-0.0234375,-0.015625,-0.0625,-0.0546875,0.1015625,0.0546875,0.0390625,-0.0078125,0.015625,-0.03125,-0.0390625,-0.0625,-0.046875,0.0546875,0.0234375,-0.03125,-0.0078125,0.0078125,-0.0546875,-0.0,-0.0234375,-0.0078125,0.0234375,-0.0390625,-0.0390625,-0.03125,0.0703125,-0.0546875,0.0625,0.0703125,-0.0625,-0.03125,-0.078125,0.015625,0.015625,0.015625,0.0390625,-0.0078125,-0.015625,-0.0390625,-0.03125,-0.0234375,0.0,-0.046875,-0.03125,-0.015625,-0.0546875,-0.046875,0.03125,0.015625,0.015625,-0.0625,0.015625,-0.0546875,-0.0234375,-0.0078125,-0.0703125,0.0078125,0.0078125,-0.0078125,-0.0078125,-0.0078125,-0.03125,0.125,-0.0625,0.0390625,-0.0078125,-0.046875,0.0390625,-0.046875,0.0625,0.1015625,-0.03125,-0.03125,-0.015625,-0.0625,0.046875,0.0,0.0234375,-0.0546875,0.0234375,-0.046875,0.0,0.0078125,0.0078125,-0.0234375,0.015625,-0.0078125,-0.0234375,-0.03125,-0.015625,-0.03125,-0.015625,0.0078125,0.0390625,-0.0234375,0.09375,0.078125,0.078125,-0.046875,-0.0390625,-0.03125,0.03125,0.0078125,-0.015625,0.0703125,0.0546875,0.015625,-0.0078125,0.203125,-0.0546875,0.0078125,-0.0078125,-0.03125,-0.0078125,-0.0078125,0.015625,0.0078125,0.0,-0.0,-0.0078125,0.0078125,-0.0078125,0.03125,-0.0546875,-0.0390625,0.0703125,-0.0078125,-0.03125,-0.0234375,-0.0234375,-0.0625,-0.0078125,0.0390625,0.0078125,0.046875,0.046875,-0.0078125,0.0625,0.0078125,-0.015625,-0.0390625,-0.0234375,-0.0703125,-0.0390625,-0.0078125,-0.03125,0.015625,0.0,-0.0625,0.015625,-0.0078125,-0.0078125,0.0,0.015625,-0.0078125,0.0,0.0078125,0.0,-0.0390625,-0.015625,-0.046875,-0.0078125,-0.03125,-0.015625,0.0390625,-0.0078125,0.015625,0.0703125,-0.0390625,0.09375,-0.046875,0.0234375,-0.078125,-0.0078125,-0.0078125,-0.0234375,0.046875,0.03125,0.0234375,0.0,-0.046875,-0.03125,-0.0234375,-0.1171875,0.0078125,0.0625,-0.0546875,-0.015625,-0.03125,0.0234375,-0.015625,-0.0703125,-0.0234375,0.0,-0.078125,0.0234375,-0.0703125,-0.0234375,0.0234375,-0.0,0.1328125,-0.015625,0.1484375,-0.0,0.0078125,0.03125,-0.03125,-0.046875,-0.046875,-0.015625,-0.015625,-0.0390625,0.046875,-0.0234375,0.015625,-0.015625,-0.0625,0.0078125,-0.015625,-0.0078125,0.0390625,-0.0078125,-0.0078125,0.0234375,-0.046875,-0.0390625,-0.03125,0.0390625,0.015625,-0.015625,-0.015625,-0.0,-0.015625,-0.046875,0.0703125,-0.0546875,0.03125,-0.046875,0.015625,0.0,-0.078125,-0.078125,0.0078125,-0.046875,0.0390625,0.015625,-0.0078125,0.0390625,0.015625,0.0,0.0078125,0.0,-0.0078125,-0.0234375,0.015625,0.0234375,-0.0078125,0.0390625,0.0,-0.015625,-0.0390625,-0.0234375,-0.0546875,0.015625,0.0078125,-0.0390625,0.015625,0.046875,0.0234375,0.046875,0.0390625,-0.0703125,-0.0078125,0.046875,-0.0390625,-0.0078125,0.03125,0.015625,-0.0546875,0.0234375,-0.046875,-0.109375,-0.0390625,-0.0546875,0.0078125,-0.0859375,-0.015625,0.0078125,-0.015625,-0.0234375,-0.0859375,0.0078125,-0.046875,0.015625,-0.0078125,0.0,-0.0078125,-0.03125,0.03125,0.0546875,-0.0703125,0.0625,0.015625,-0.0,0.0703125,0.0234375,-0.0703125,-0.0390625,-0.0,0.0,-0.03125,0.078125,-0.0625,0.0,0.046875,-0.125,0.0546875,0.0078125,-0.0,-0.0625,0.015625,0.0078125,-0.0,-0.046875,-0.03125,-0.0,0.015625,-0.078125,-0.03125,0.0625,-0.03125,0.1171875,0.0,-0.0390625,0.0546875,-0.0546875,-0.0390625,-0.03125,0.03125,0.0078125,0.015625,0.0078125,-0.015625,-0.0546875,-0.0703125,-0.03125,-0.046875,0.046875,-0.1171875,0.0,0.0859375,-0.0390625,0.0859375,-0.046875,-0.1015625,0.03125,-0.0546875,-0.0546875,-0.0078125,-0.015625,-0.0625,-0.0546875,0.0390625,0.1171875,0.078125,0.0546875,-0.03125,0.0234375,-0.0625,-0.0390625,0.015625,-0.03125,0.0859375,0.109375,-0.0078125,-0.0234375,0.0625,-0.046875,0.03125,0.015625,-0.0625,-0.0,-0.0234375,0.0546875,-0.0625,0.015625,0.0546875,0.03125,0.0625,0.0234375,-0.046875,0.015625,-0.0078125,-0.0859375,-0.015625,-0.0078125,0.015625,0.0859375,0.03125,-0.0078125,0.0234375,0.015625,-0.0078125,-0.0078125,0.0,0.015625,-0.015625,-0.0078125,-0.0078125,-0.015625,-0.03125,-0.0234375,-0.0390625,0.0625,-0.078125,0.046875,0.0390625,-0.0078125,0.046875,-0.0078125,-0.0078125,0.0546875,-0.0078125,-0.0625,-0.0234375,0.0703125,-0.0390625,0.0390625,-0.0390625,0.0078125,0.0,-0.03125,0.0859375,0.0546875,-0.015625,-0.015625,-0.0625,0.0,-0.0078125,0.0,0.0078125,-0.0078125,-0.0078125,0.0078125,0.0078125,0.0078125,-0.015625,-0.0234375,-0.0078125,0.0546875,0.03125,-0.015625,-0.0,0.0390625,-0.0625,-0.015625,-0.0234375,-0.0234375,0.1015625,-0.015625,0.15625,0.0546875,-0.0625,0.0234375,0.0234375,0.0,0.0078125,-0.0703125,-0.03125,-0.0,-0.046875,-0.0234375,0.046875,0.0078125,0.03125,0.0078125,0.015625,0.0,0.0078125,-0.0078125,-0.0078125,0.015625,-0.0234375,-0.0859375,-0.0234375,-0.0,-0.09375,0.046875,0.015625,0.015625,-0.0,-0.0234375,-0.0390625,-0.0078125,0.0,-0.0390625,-0.0234375,-0.0,-0.015625,0.015625,0.0,-0.03125,-0.03125,0.0625,-0.0078125,0.0546875,0.0078125,-0.0,0.0390625,0.015625,0.0078125,-0.0078125,0.03125,0.03125,-0.046875,-0.03125,0.0,-0.0234375,-0.03125,-0.0234375,0.0078125,-0.0390625,0.03125,-0.0390625,0.046875,-0.046875,0.0078125,0.0078125,0.015625,-0.0078125,-0.0234375,0.1015625,0.0859375,-0.0,0.0390625,-0.0234375,-0.0,-0.0078125,0.0,-0.0078125,-0.015625,-0.015625,0.0078125,-0.0,0.0,-0.015625,0.0078125,-0.046875,0.0234375,-0.0546875,-0.0625,0.0078125,-0.03125,-0.0078125,-0.03125,0.0234375,0.03125,-0.03125,0.0078125,-0.015625,-0.0078125,-0.03125,-0.0,-0.0,-0.0,0.046875,-0.03125,0.0546875,-0.0234375,-0.0390625,-0.1328125,-0.0390625,-0.015625,-0.0546875,0.0234375,0.0234375,0.078125,0.046875,0.015625,-0.0078125,-0.0078125,-0.0078125,-0.03125,0.1015625,0.046875,0.0390625,0.0078125,-0.0390625,-0.078125,-0.0625,-0.0234375,-0.03125,-0.0390625,0.0546875,-0.0078125,0.0078125,-0.0234375,-0.03125,0.0703125,-0.0390625,-0.015625,-0.0078125,-0.09375,0.0234375,-0.0546875,0.046875,0.0078125,-0.0390625,-0.0234375,-0.0078125,-0.015625,-0.046875,-0.046875,-0.046875,-0.015625,-0.0234375,0.015625,-0.0078125,0.015625,0.0234375,-0.0546875,-0.1328125,-0.0625,-0.078125,-0.0546875,-0.0625,-0.0234375,-0.03125,0.015625,0.0546875,0.0390625,0.015625,0.0078125,0.046875,0.0546875,-0.046875,0.0546875,-0.015625,0.0390625,-0.015625,-0.078125,-0.03125,-0.0703125,-0.1171875,0.015625,-0.0234375,0.0078125,-0.0703125,0.0546875,0.0,-0.0234375,0.0234375,-0.0625,-0.03125,0.09375,-0.0078125,-0.0234375,-0.1015625,-0.0,0.0234375,-0.03125,-0.015625,0.015625,-0.0234375,-0.0390625,0.03125,0.0390625,0.0859375,-0.015625,0.03125,-0.0078125,-0.0234375,0.03125,-0.015625,-0.078125,-0.046875,-0.03125,-0.0,-0.03125,-0.0234375,0.0390625,0.0078125,0.03125,0.0,-0.0078125,0.09375,0.0078125,-0.0,-0.046875,-0.015625,0.0078125,0.0,0.0078125,-0.0078125,-0.015625,-0.0,-0.0,-0.0078125,-0.015625,0.03125,0.0078125,-0.0234375,0.0,0.015625,0.0078125,0.0234375,-0.0078125,0.046875,-0.0546875,-0.03125,0.0546875,0.0078125,-0.0234375,0.015625,-0.015625,0.0,0.03125,0.1640625,-0.0390625,0.0546875,0.0078125,-0.078125,-0.0703125,-0.0234375,-0.015625,-0.0,-0.0078125,0.015625,0.0078125,-0.0078125,0.015625,-0.0,0.0078125,0.015625,0.0390625,0.0625,0.015625,-0.015625,-0.0625,-0.1015625,-0.03125,0.03125,0.015625,0.0234375,0.078125,-0.0078125,-0.015625,0.015625,0.0390625,0.0390625,-0.0078125,-0.03125,-0.0703125,0.125,0.015625,0.0,-0.03125,-0.0390625,0.0078125,-0.03125,0.0390625,0.0234375,0.0078125,-0.015625,0.015625,0.03125,0.03125,-0.0234375,0.0078125,-0.0078125,-0.0390625,0.015625,0.0,0.0703125,0.0703125,-0.03125,-0.0234375,-0.03125,-0.0078125,0.0390625,0.0078125,-0.046875,-0.03125,-0.03125,-0.0546875,-0.0390625,-0.03125,-0.0234375,-0.0078125,0.0078125,0.0078125,-0.0078125,-0.0,0.0,0.0,0.0078125,-0.015625,-0.0234375,0.0234375,0.0234375,-0.046875,-0.078125,-0.015625,0.015625,0.015625,0.0546875,-0.03125,0.015625,0.0546875,0.0703125,-0.1015625,-0.03125,0.046875,-0.0078125,0.015625,-0.0390625,0.03125,0.046875,-0.1015625,-0.078125,0.015625,0.0234375,0.03125,-0.0,0.0078125,-0.0078125,0.0,-0.0,0.0078125,-0.0,-0.0,-0.0,-0.015625,0.0234375,-0.046875,0.0234375,0.0078125,-0.0,-0.0234375,-0.03125,-0.0390625,-0.03125,-0.0625,-0.0546875,-0.03125,-0.0234375,0.03125,0.0234375,-0.0546875,0.015625,-0.046875,-0.0390625,0.09375,-0.0234375,0.0078125,0.0703125,-0.0859375,0.0390625,0.0234375,-0.015625,-0.0,-0.03125,-0.0234375,-0.0859375,-0.03125,-0.078125,-0.0078125,0.0234375,0.0078125,0.078125,0.0,0.0390625,-0.0078125,-0.0390625,0.015625,-0.0078125,-0.0234375,0.0234375,0.0234375,0.09375,0.0234375,-0.03125,0.0390625,-0.015625,-0.015625,0.03125,-0.015625,-0.0078125,-0.0546875,-0.046875,0.0234375,-0.0,0.0,-0.0390625,-0.0078125,-0.03125,0.0703125,-0.0390625,0.03125,0.015625,0.0,-0.078125,-0.0625,-0.0234375,0.0,0.015625,0.0703125,0.0,-0.03125,-0.0625,0.0,-0.078125,0.0,-0.046875,-0.046875,0.0546875,0.0546875,-0.0546875,0.0625,0.0,-0.0078125,-0.0390625,0.0078125,0.0078125,0.0078125,0.0078125,-0.0703125,-0.125,-0.0234375,-0.0234375,-0.0234375,0.0703125,-0.0078125,-0.0,-0.0703125,0.125,-0.0234375,0.0078125,-0.0234375,0.0234375,0.0,-0.0546875,0.0078125,-0.046875,-0.0078125,-0.0390625,0.046875,-0.0546875,0.03125,-0.0078125,-0.0625,0.125,0.03125,-0.0234375,0.03125,0.015625,0.0078125,0.015625,-0.0234375,0.0078125,-0.0234375,0.0078125,-0.046875,0.015625,0.0546875,-0.015625,-0.0546875,-0.0546875,-0.03125,-0.03125,-0.03125,-0.03125,0.0546875,-0.0078125,-0.0390625,-0.0234375,-0.015625,0.0,-0.015625,-0.0078125,-0.0078125,0.0078125,0.0,0.015625,0.015625,-0.0,-0.015625,0.0078125,-0.0234375,0.0078125,-0.0390625,-0.0390625,-0.046875,-0.0390625,0.0078125,0.03125,-0.03125,0.0390625,-0.0,0.0078125,-0.0078125,-0.03125,0.0078125,-0.015625,0.0625,0.078125,-0.0625,-0.0703125,-0.0390625,-0.0234375,-0.0,-0.03125,0.0,0.0078125,-0.0,-0.0078125,-0.0078125,0.0,0.0078125,0.0,0.0,0.0078125,0.0234375,0.0078125,0.0546875,-0.0234375,0.0,-0.0234375,0.0546875,-0.03125,-0.0390625,0.03125,-0.0078125,-0.0078125,-0.0703125,-0.0078125,-0.0390625,0.0078125,0.0234375,-0.0,-0.0390625,-0.0078125,0.0078125,0.0390625,0.09375,-0.0546875,-0.0,-0.015625,-0.03125,-0.0078125,-0.0390625,-0.03125,0.078125,0.015625,0.0078125,-0.015625,0.0078125,0.0390625,-0.0546875,-0.0234375,0.03125,-0.0703125,-0.0234375,0.0078125,-0.0234375,0.0,-0.015625,-0.0,0.015625,0.0078125,-0.015625,0.0078125,0.0,0.015625,0.0234375,-0.015625,-0.0078125,0.0,0.015625,0.015625,0.0078125,-0.0234375,-0.0,0.0078125,0.0078125,0.0078125,-0.0078125,-0.0,0.0390625,0.0,-0.03125,-0.0,-0.046875,-0.0,-0.0390625,0.015625,-0.0078125,-0.0078125,0.109375,-0.0,-0.046875,-0.0234375,-0.0390625,-0.015625,-0.015625,-0.015625,0.0078125,0.03125,-0.03125,0.015625,-0.0078125,-0.0078125,-0.0,0.015625,0.0,-0.015625,-0.015625,-0.015625,0.0078125,0.0078125,0.0078125,0.015625,-0.0234375,0.03125,0.0,-0.0,-0.03125,-0.0234375,0.0078125,-0.0078125,0.0546875,0.0078125,-0.0,0.015625,-0.0546875,-0.015625,-0.0078125,-0.0,0.0078125,0.0078125,0.03125,-0.0078125,0.0234375,0.0546875,0.03125,-0.0390625,-0.015625,-0.0234375,0.0703125,0.0,-0.03125,-0.0625,-0.0703125,-0.046875,0.0625,-0.0,-0.0234375,-0.0234375,-0.0234375,0.0,0.0234375,-0.046875,-0.03125,-0.0390625,-0.0234375,0.0234375,-0.015625,-0.0078125,-0.03125,-0.0234375,0.0078125,-0.0078125,-0.015625,0.0078125,-0.0,0.046875,0.015625,-0.0,0.078125,-0.03125,-0.046875,0.0078125,-0.015625,0.0234375,-0.0390625,-0.0,-0.0078125,0.015625,0.0078125,-0.0078125,-0.03125,-0.0078125,-0.015625,-0.0078125,0.046875,0.015625,0.0625,0.0078125,-0.0,0.0234375,-0.015625,-0.0,-0.046875,-0.046875,0.0,-0.09375,-0.0859375,-0.03125,-0.0390625,0.0078125,0.0,0.09375,-0.046875,-0.046875,0.1171875,-0.0546875,0.0234375,-0.0234375,-0.046875,-0.015625,0.0078125,0.078125,0.015625,-0.09375,-0.0078125,-0.015625,-0.0,0.0078125,0.015625,-0.015625,-0.03125,-0.0078125,-0.0234375,0.015625,0.0234375,-0.03125,-0.0703125,0.0625,-0.03125,0.0859375,-0.0078125,-0.0078125,0.0234375,0.0,0.0390625,0.0078125,0.015625,0.015625,-0.0078125,-0.0,0.078125,-0.1015625,0.015625,0.0,0.0,0.0390625,0.0546875,-0.0625,0.0078125,-0.0625,-0.015625,0.0,-0.0234375,-0.0625,0.125,0.0078125,-0.0078125,-0.0078125,0.0234375,-0.0,0.0,-0.0078125,0.0078125,0.015625,-0.0234375,-0.0234375,0.0078125,0.0078125,-0.046875,0.140625,0.0234375,-0.046875,-0.015625,-0.0078125,0.0390625,0.0,-0.015625,-0.0546875,0.078125,0.0234375,0.015625,-0.0078125,0.03125,0.0859375,-0.015625,-0.0234375,-0.0625,-0.03125,-0.0390625,0.03125,-0.015625,0.015625,-0.0078125,0.0078125,0.0078125,0.0078125,0.015625,-0.015625,-0.0078125,0.0,0.0234375,0.0078125,-0.0390625,0.0,0.0390625,-0.03125,0.03125,-0.0625,0.0078125,-0.0234375,-0.0234375,0.03125,0.0,-0.0234375,0.0078125,0.015625,-0.0390625,0.015625,0.0546875,0.0,-0.0546875,-0.0859375,-0.046875,-0.046875,0.0,-0.046875,0.03125,-0.046875,-0.046875,-0.0390625,0.0078125,-0.015625,-0.0390625,0.03125,-0.03125,-0.0078125,0.046875,-0.046875,-0.0078125,0.0078125,-0.03125,-0.015625,-0.0859375,0.03125,0.046875,-0.0078125,0.0625,0.0078125,0.0390625,0.015625,-0.015625,0.0078125,0.0078125,0.015625,-0.0,-0.015625,-0.015625,0.0078125,0.03125,0.0078125,-0.015625,0.015625,-0.015625,0.0234375,0.0078125,0.015625,-0.0234375,-0.0078125,-0.0234375,-0.03125,-0.015625,-0.0234375,0.1171875,-0.0625,-0.03125,-0.0234375,-0.0234375,-0.03125,-0.046875,-0.015625,0.0546875,0.0390625,0.0078125,-0.0234375,-0.0234375,-0.0,0.03125,-0.0390625,0.0,-0.0,-0.015625,-0.0078125,0.0078125,-0.0078125,0.0234375,0.0234375,-0.0078125,-0.0,-0.0078125,-0.015625,-0.03125,-0.015625,0.03125,-0.0078125,-0.0,0.0234375,0.0,0.015625,-0.0078125,-0.0234375,-0.0,-0.03125,0.0078125,-0.0078125,-0.046875,0.015625,-0.0078125,-0.0078125,-0.0390625,-0.0,0.0078125,-0.015625,0.0,-0.03125,0.0390625,-0.015625,0.03125,-0.0546875,0.015625,-0.0234375,0.0,0.0078125,-0.0390625,0.046875,0.0625,0.0234375,0.0078125,-0.0234375,0.0390625,0.03125,-0.046875,-0.0625,-0.0234375,-0.046875,-0.0625,-0.046875,-0.0,0.0703125,0.015625,0.046875,0.046875,-0.0234375,-0.015625,0.0625,-0.0,0.078125,-0.015625,-0.1171875,-0.0859375,-0.0078125,0.0234375,-0.0390625,-0.0390625,-0.0,-0.0234375,0.0625,-0.046875,-0.0,-0.0390625,0.015625,0.0234375,0.03125,0.0078125,-0.015625,0.0703125,0.0,-0.0078125,0.0546875,0.0390625,-0.0390625,-0.0234375,0.0546875,0.0703125,-0.0703125,0.078125,0.0546875,-0.015625,-0.015625,-0.0546875,-0.03125,-0.0078125,0.0078125,-0.046875,-0.0625,-0.0078125,0.015625,0.03125,-0.03125,0.0078125,-0.03125,-0.0078125,-0.03125,0.015625,-0.0546875,-0.0078125,0.078125,0.0234375,-0.0234375,0.0234375,-0.0078125,0.0625,0.0390625,-0.03125,0.03125,-0.015625,-0.0625,0.015625,-0.0546875,-0.0390625,0.1015625,0.0390625,-0.0546875,0.046875,0.0390625,0.0078125,0.0078125,0.015625,-0.0078125,-0.0078125,-0.03125,-0.078125,-0.0390625,-0.0078125,-0.046875,0.015625,0.0,0.0078125,-0.0703125,0.0546875,-0.0078125,0.0546875,-0.015625,0.0390625,0.0,0.0078125,-0.0078125,0.0,0.015625,-0.0,-0.0,-0.0,0.0,-0.015625,-0.0390625,0.046875,0.0078125,-0.046875,0.0546875,-0.0234375,-0.1328125,-0.0703125,-0.0078125,-0.0234375,-0.0,0.0625,-0.03125,0.0625,-0.078125,-0.0078125,-0.0390625,0.0390625,0.0546875,0.03125,-0.09375,-0.0390625,-0.03125,0.015625,0.046875,0.140625,0.0078125,0.015625,0.0,-0.0,0.0,0.0,-0.0078125,-0.015625,-0.0,-0.03125,0.0546875,0.03125,-0.015625,-0.0234375,0.0625,0.0703125,-0.015625,-0.0625,-0.03125,0.0078125,-0.015625,0.0234375,-0.046875,-0.015625,0.046875,-0.046875,0.0546875,0.0078125,-0.0625,-0.03125,-0.0078125,-0.0703125,-0.0078125,-0.0078125,-0.015625,0.015625,0.0078125,-0.03125,-0.0,-0.0078125,0.0234375,0.0,0.0390625,-0.109375,-0.03125,-0.0078125,-0.0078125,-0.0859375,0.046875,0.0625,-0.0390625,-0.078125,-0.0703125,-0.0390625,-0.0078125,0.0078125,0.0,-0.0390625,0.0078125,0.0078125,0.0546875,0.03125,-0.015625,-0.0390625,0.015625,0.0078125,0.0078125,-0.0390625,0.03125,0.0078125,-0.0546875,-0.015625,0.0234375,0.0078125,0.0,-0.0078125,-0.0390625,0.0546875,0.015625,0.0625,0.015625,-0.0234375,0.015625,-0.0078125,0.0078125,-0.0234375,-0.03125,0.0859375,-0.0390625,0.0703125,0.03125,0.0390625,0.0390625,-0.0234375,-0.0859375,-0.078125,0.046875,-0.0546875,0.015625,-0.0,-0.0078125,-0.0078125,-0.0,0.0078125,0.0078125,-0.0,-0.015625,0.0078125,-0.0,-0.0078125,0.0234375,0.03125,-0.0,0.0078125,0.0,-0.046875,0.0078125,-0.0546875,-0.015625,-0.046875,0.0078125,-0.0546875,0.1015625,-0.1328125,-0.015625,0.0234375,-0.0,0.015625,0.0078125,-0.015625,-0.0234375,0.03125,0.109375,0.046875,-0.0234375,-0.015625,0.0234375,-0.0078125,-0.0546875,-0.0234375,0.0078125,-0.0546875,0.0390625,0.0390625,-0.0,-0.0078125,-0.0390625,-0.1015625,-0.046875,-0.0078125,0.1015625,-0.015625,-0.0078125,0.0625,-0.0390625,0.0,-0.0625,0.0234375,-0.015625,-0.0,0.046875,-0.0703125,-0.015625,-0.0546875,-0.0546875,0.0,0.03125,0.0234375,-0.15625,0.078125,-0.03125,0.0546875,0.015625,-0.03125,-0.0234375,0.0546875,-0.0546875,-0.0703125,0.0234375,-0.0625,0.0390625,-0.0234375,0.0078125,0.046875,-0.0078125,-0.1015625,0.015625,0.015625,-0.0,0.03125,0.03125,0.0078125,0.0390625,-0.09375,0.0390625,0.046875,-0.0546875,-0.015625,-0.015625,-0.0390625,-0.03125,0.0390625,-0.1484375,0.0546875,0.0546875,-0.0703125,0.078125,-0.046875,0.0078125,-0.046875,-0.0390625,0.0703125,0.109375,-0.0234375,-0.0234375,0.09375,-0.0234375,-0.0390625,-0.03125,0.125,-0.03125,0.03125,-0.0390625,-0.015625,-0.125,-0.0390625,-0.0078125,-0.015625,0.046875,0.1015625,-0.0390625,-0.0546875,0.0546875,-0.0625,-0.015625,-0.0,0.0390625,0.0078125,0.0625,-0.03125,-0.0234375,0.0078125,-0.0234375,0.0234375,-0.015625,-0.0078125,-0.0,0.078125,-0.0234375,-0.0234375,0.078125,0.03125,0.0,-0.0078125,-0.015625,0.0078125,-0.0078125,0.0078125,-0.0078125,0.0078125,0.015625,0.0078125,-0.0234375,0.0078125,0.015625,-0.0546875,-0.0625,0.0234375,-0.0234375,0.0859375,0.0,-0.0234375,0.015625,0.0078125,0.03125,-0.0078125,-0.03125,-0.0078125,-0.0234375,-0.015625,0.0078125,-0.015625,-0.0078125,-0.0234375,-0.015625,-0.0078125,-0.0078125,0.0703125,0.0078125,-0.0,0.0,-0.0,0.0,-0.0,0.0078125,0.0078125,-0.015625,-0.0234375,-0.03125,-0.0078125,-0.0234375,0.03125,0.0234375,-0.0,-0.0078125,-0.0078125,0.0,-0.0,-0.046875,-0.0234375,-0.046875,0.0390625,-0.0390625,0.0234375,0.09375,0.0,0.046875,0.0234375,-0.0078125,-0.0234375,-0.046875,-0.0234375,-0.1015625,0.0390625,0.015625,-0.03125,-0.0234375,-0.0078125,-0.0625,-0.0390625,-0.0078125,0.0,0.015625,0.0078125,-0.0234375,-0.0234375,-0.0234375,0.03125,0.046875,-0.0078125,-0.0078125,-0.0,-0.0,-0.0,-0.0234375,-0.03125,0.0078125,0.0,0.0,0.0234375,0.0625,0.015625,0.0078125,0.0,0.015625,-0.0,0.0234375,0.0078125,0.0078125,0.0078125,0.0078125,0.0078125,0.0078125,0.0078125,-0.0078125,-0.015625,0.0390625,-0.0390625,-0.0546875,-0.0,0.015625,-0.0234375,-0.015625,0.0078125,0.0078125,-0.015625,0.0859375,-0.0390625,-0.015625,-0.015625,-0.0078125,-0.0234375,-0.0390625,0.0078125,0.0390625,-0.015625,-0.03125,-0.0078125,0.0,-0.0,0.0078125,-0.0078125,0.0078125,0.0078125,0.0078125,0.0234375,0.015625,-0.0078125,-0.0234375,-0.015625,-0.015625,-0.0078125,0.0078125,-0.0390625,0.0078125,-0.015625,-0.015625,0.0234375,-0.015625,-0.0234375,-0.0546875,0.0,-0.0078125,-0.0234375,-0.0078125,-0.0390625,-0.03125,-0.03125,-0.0234375,0.0234375,-0.0234375,-0.0234375,0.078125,0.0,-0.0078125,-0.015625,-0.0390625,-0.0859375,-0.046875,0.0234375,0.0078125,-0.046875,0.015625,-0.015625,-0.0390625,-0.015625,0.03125,0.0,0.03125,0.03125,0.03125,-0.0,0.0234375,0.015625,0.015625,-0.0234375,-0.03125,0.0234375,0.03125,0.0390625,-0.015625,-0.0078125,-0.0234375,-0.015625,-0.0546875,0.0,-0.0,-0.0703125,0.0625,0.0078125,-0.0078125,0.015625,-0.0078125,-0.046875,-0.03125,-0.015625,-0.015625,0.0078125,-0.015625,0.015625,-0.0,0.0078125,0.0234375,-0.0234375,-0.0078125,-0.0,-0.0,-0.0,-0.03125,-0.0234375,-0.0234375,0.0,0.1015625,0.0390625,-0.03125,0.015625,-0.015625,0.015625,-0.0234375,-0.0234375,0.015625,-0.0625,0.015625,0.0546875,-0.0703125,0.0078125,0.0,-0.0078125,-0.0078125,-0.0078125,-0.015625,-0.03125,-0.0234375,-0.03125,-0.015625,-0.0,-0.0,0.015625,-0.015625,0.03125,0.015625,-0.0,-0.0625,-0.015625,-0.0,-0.015625,0.03125,-0.03125,0.0078125,0.0,-0.046875,0.0,0.0078125,-0.0078125,-0.03125,-0.046875,0.046875,-0.0,-0.0078125,-0.015625,0.0390625,-0.0078125,-0.046875,-0.0703125,0.0390625,-0.046875,0.046875,0.1015625,0.0234375,-0.0078125,-0.0078125,-0.0078125,0.0078125,-0.015625,-0.0078125,-0.0234375,0.0078125,0.0,-0.0078125,0.03125,0.0,-0.03125,-0.09375,-0.1015625,0.015625,-0.0078125,-0.03125,-0.0078125,0.015625,-0.015625,-0.0703125,0.0078125,-0.0390625,-0.0390625,-0.0078125,-0.046875,0.0078125,-0.046875,0.0078125,0.0546875,-0.0078125,-0.0078125,-0.046875,-0.0234375,0.09375,-0.125,-0.0078125,-0.015625,0.0078125,0.0078125,0.0078125,0.015625,0.0078125,-0.0,0.0078125,-0.0546875,-0.0390625,0.015625,0.0078125,-0.03125,-0.0390625,0.03125,0.0859375,-0.078125,0.1484375,0.078125,-0.046875,0.046875,-0.0625,-0.0390625,0.0625,-0.015625,-0.015625,-0.0234375,-0.0078125,-0.09375,-0.0078125,-0.0546875,-0.0078125,0.078125,0.078125,-0.0703125,-0.0078125,0.0078125,-0.0,-0.0078125,-0.0078125,0.0078125,-0.0390625,0.0078125,0.0078125,-0.0390625,0.0078125,0.015625,0.015625,0.03125,0.1015625,-0.046875,-0.0390625,-0.0078125,-0.03125,-0.0625,0.0390625,0.0625,0.0625,-0.0234375,-0.0,-0.0625,0.015625,-0.0234375,0.09375,-0.015625,-0.0234375,0.0,-0.0,-0.046875,0.0078125,0.0078125,-0.046875,-0.0234375,-0.046875,0.0546875,0.0234375,-0.0390625,-0.046875,0.0234375,0.015625,-0.015625,0.015625,0.0390625,0.078125,0.015625,0.046875,-0.0390625,-0.0390625,-0.0234375,0.0546875,-0.0703125,0.109375,0.0078125,-0.140625,-0.0078125,0.0390625,0.0546875,-0.0234375,-0.0078125,-0.015625,-0.03125,-0.015625,-0.0234375,-0.0234375,0.0078125,0.0,-0.0078125,-0.0078125,-0.0078125,-0.0390625,0.015625,0.0703125,-0.046875,-0.0546875,-0.0078125,0.0546875,0.03125,-0.015625,-0.0625,-0.0859375,-0.0078125,-0.0078125,-0.0,-0.0234375,0.046875,-0.015625,-0.015625,0.0390625,-0.0234375,-0.03125,-0.0546875,0.0625,0.125,-0.0625,-0.0078125,0.0078125,0.046875,-0.1171875,-0.046875,-0.015625,-0.046875,-0.0546875,0.0546875,-0.0625,-0.0546875,-0.0390625,-0.0390625,-0.0234375,0.0078125,0.0390625,-0.0390625,-0.0234375,0.0625,-0.0703125,0.03125,-0.0625,-0.0078125,0.0546875,0.0234375,0.0390625,0.0,0.078125,0.0,0.0078125,-0.0234375,-0.0078125,0.0390625,-0.078125,-0.078125,0.140625,-0.09375,-0.0703125,0.0703125,-0.0546875,0.0546875,0.0703125,-0.1015625,-0.0703125,0.046875,0.0390625,0.0078125,0.046875,-0.015625,-0.0234375,0.0625,0.0234375,0.0390625,0.0,-0.0859375,-0.0390625,-0.0078125,0.0,0.03125,0.0,0.0,0.1328125,-0.015625,0.0859375,0.03125,0.015625,-0.0078125,-0.015625,-0.0390625,-0.015625,-0.0390625,0.0,-0.0234375,-0.09375,0.0546875,0.015625,-0.0078125,-0.109375,-0.0390625,-0.1171875,-0.015625,0.0703125,0.1328125,-0.0546875,-0.03125,0.0546875,-0.1015625,-0.078125,0.03125,0.03125,0.0625,-0.0390625,0.125,0.0078125,-0.03125,-0.015625,0.0078125,0.015625,0.0234375,0.046875,0.015625,-0.0390625,0.0078125,-0.1640625,-0.0625,-0.0234375,-0.046875,-0.0234375,-0.015625,-0.03125,-0.0546875,-0.078125,-0.015625,0.0,0.078125,0.0703125,0.0390625,-0.0078125,-0.015625,0.015625,-0.0078125,0.0078125,-0.0,0.015625,-0.0078125,-0.0,0.0078125,-0.0234375,-0.03125,-0.0078125,-0.078125,0.0703125,0.0625,-0.0390625,-0.0390625,0.0625,0.0390625,-0.0859375,-0.0234375,-0.0390625,-0.0546875,0.015625,0.03125,-0.0390625,-0.0,-0.015625,0.046875,0.03125,-0.03125,0.078125,-0.03125,-0.0390625,0.0078125,-0.0078125,0.0078125,0.0078125,-0.0078125,0.0,0.0078125,0.015625,0.0078125,-0.0078125,0.0078125,-0.0234375,0.0234375,-0.0078125,0.0078125,0.015625,0.0234375,0.0,-0.0,0.0390625,-0.1640625,-0.015625,0.0078125,-0.0078125,-0.0625,-0.0078125,0.0234375,0.015625,-0.046875,-0.03125,-0.0234375,0.0,-0.0703125,0.0546875,-0.0234375,-0.0234375,-0.0234375,-0.0390625,-0.0078125,0.1171875,0.0078125,-0.015625,0.0,0.0234375,-0.0234375,0.0078125,0.015625,-0.0,-0.0234375,-0.0390625,0.015625,-0.0703125,-0.03125,-0.0625,-0.03125,-0.03125,-0.015625,-0.0078125,0.046875,0.03125,-0.015625,0.0078125,-0.0234375,-0.0234375,-0.0,0.0234375,-0.03125,-0.015625,-0.0546875,0.0078125,0.0234375,-0.0078125,0.0,-0.0234375,0.0234375,-0.0234375,0.0703125,-0.0625,-0.0078125,0.0234375,-0.0234375,-0.0234375,-0.03125,0.03125,0.0234375,0.0234375,-0.0078125,-0.0234375,-0.03125,0.0078125,-0.0390625,0.03125,0.109375,0.0390625,-0.03125,-0.046875,0.0546875,0.015625,-0.0859375,-0.0078125,0.0,0.015625,0.0078125,-0.0234375,0.0234375,-0.0,0.0078125,0.015625,-0.0234375,-0.0234375,-0.0625,-0.03125,-0.0078125,-0.0078125,0.0078125,-0.0078125,0.03125,-0.0,0.0546875,-0.015625,0.0,0.078125,-0.03125,0.0,0.0,0.015625,-0.0078125,-0.0078125,-0.0703125,0.046875,0.0234375,-0.09375,-0.0234375,-0.015625,-0.0625,-0.0625,0.0078125,-0.1171875,0.0546875,0.0625,0.0859375,0.03125,-0.03125,-0.015625,-0.03125,-0.0546875,-0.046875,0.0390625,-0.0234375,-0.03125,0.0078125,-0.0390625,-0.0,-0.0234375,-0.0390625,0.0859375,-0.0703125,-0.015625,-0.0234375,0.0703125,-0.015625,0.015625,-0.0234375,0.0703125,0.1640625,-0.078125,-0.046875,-0.0390625,0.0,-0.0,0.0234375,-0.0546875,0.015625,-0.0546875,-0.0546875,0.0,0.0,0.015625,0.0078125,-0.0078125,-0.0078125,-0.015625,0.0078125,-0.03125,0.015625,-0.0625,-0.0078125,-0.0703125,-0.015625,0.0078125,-0.0078125,-0.0546875,-0.03125,0.046875,0.0703125,0.0,0.0078125,-0.0703125,-0.015625,-0.1484375,-0.0234375,-0.09375,-0.0234375,0.0390625,0.015625,0.0546875,-0.0625,-0.0,0.0,-0.0390625,0.0625,0.0234375,0.0234375,-0.0078125,-0.0234375,-0.0625,0.015625,0.0625,0.1171875,-0.015625,0.0234375,-0.015625,-0.0390625,-0.0234375,-0.0078125,-0.015625,-0.1015625,0.0234375,0.0078125,0.015625,0.0390625,0.0546875,0.03125,0.0078125,0.0234375,0.0078125,0.0078125,-0.09375,-0.03125,-0.0859375,-0.046875,0.0078125,0.0859375,0.015625,0.015625,0.0625,0.03125,0.09375,-0.03125,0.015625,0.0390625,-0.015625,-0.0234375,-0.015625,-0.015625,0.0078125,0.015625,0.0078125,-0.0078125,0.015625,0.0078125,-0.015625,-0.0390625,-0.015625,0.1328125,-0.03125,-0.0078125,-0.0234375,0.0703125,0.015625,-0.0078125,-0.0078125,0.015625,0.0,0.03125,0.0234375,-0.03125,0.03125,-0.0234375,0.0078125,-0.0625,-0.015625,-0.0234375,-0.0390625,-0.0390625,-0.03125,0.03125,-0.015625,-0.0234375,-0.0078125,-0.0078125,-0.015625,-0.015625,0.0078125,0.0078125,-0.0,-0.015625,0.0078125,-0.0546875,-0.0625,-0.015625,-0.0078125,0.0390625,-0.015625,-0.109375,-0.0078125,-0.0234375,-0.125,0.0859375,-0.0390625,0.046875,-0.0703125,-0.03125,0.1484375,0.0234375,-0.0390625,-0.0859375,-0.0234375,-0.015625,0.03125,-0.015625,-0.0078125,0.1015625,-0.078125,-0.0390625,0.0390625,0.1015625,0.0078125,-0.03125,-0.0,-0.0078125,-0.046875,-0.015625,0.0234375,-0.0703125,-0.046875,-0.03125,-0.0234375,0.0390625,-0.0234375,-0.046875,-0.0625,-0.03125,-0.046875,0.0078125,-0.0,-0.0,-0.0,-0.0390625,0.09375,-0.09375,-0.0078125,-0.03125,0.0234375,0.0,-0.0390625,-0.015625,0.015625,0.0078125,0.0078125,-0.015625,0.03125,-0.0234375,-0.015625,0.0390625,-0.0390625,0.015625,-0.015625,-0.015625,-0.015625,0.0625,0.171875,-0.0,-0.125,-0.0859375,-0.046875,-0.03125,0.0,-0.0390625,-0.0625,0.0078125,-0.046875,0.0625,0.0234375,0.0,-0.0234375,-0.0234375,-0.015625,0.0078125,0.0078125,-0.0078125,-0.0,-0.03125,-0.0078125,0.015625,0.0078125,-0.0,-0.015625,-0.015625,0.0234375,-0.046875,-0.0390625,0.0234375,0.0546875,0.0078125,0.0,0.0546875,-0.0390625,0.0,0.0234375,-0.0078125,-0.0390625,0.0234375,0.0078125,-0.0234375,-0.0078125,0.046875,-0.0390625,-0.078125,-0.0234375,-0.03125,0.1484375,-0.0234375,-0.0234375,0.0625,-0.09375,-0.0390625,-0.078125,0.09375,-0.0078125,-0.03125,-0.0390625,0.0078125,-0.09375,0.0,0.0234375,-0.1171875,0.046875,0.046875,0.0859375,-0.0234375,-0.0546875,0.015625,-0.046875,0.0234375,0.0546875,-0.09375,-0.03125,0.0703125,-0.015625,-0.0546875,0.0703125,-0.0,0.03125,-0.0078125,-0.125,-0.0078125,-0.015625,-0.046875,-0.0703125,-0.0625,-0.015625,-0.0078125,-0.1015625,0.046875,-0.0078125,0.1015625,0.0234375,0.015625,0.0,-0.015625,-0.0,-0.0078125,-0.0546875,-0.015625,0.1171875,-0.0078125,-0.0234375,-0.0859375,0.03125,0.046875,0.0390625,-0.0390625,-0.0390625,0.03125,-0.078125,-0.046875,0.0390625,0.0,-0.03125,0.0625,0.046875,-0.0078125,-0.0234375,-0.0625,-0.0390625,-0.0546875,0.0078125,0.0859375,-0.0625,0.0625,-0.0625,-0.0234375,-0.015625,0.0078125,-0.03125,0.0234375,0.03125,0.0234375,-0.171875,-0.0234375,-0.03125,0.1328125,-0.046875,-0.015625,-0.078125,-0.0625,0.0703125,-0.0703125,-0.0390625,0.03125,0.0234375,-0.03125,0.015625,0.0,0.0546875,0.0,-0.0703125,0.0078125,0.0390625,-0.046875,-0.046875,-0.0078125,0.046875,-0.0546875,-0.0859375,-0.0625,0.015625,0.0234375,-0.03125,-0.03125,-0.015625,-0.015625,0.015625,0.0078125,-0.0078125,-0.0078125,0.0234375,0.0,0.0,0.0,0.015625,-0.0390625,0.0078125,0.0,-0.0078125,0.0234375,-0.03125,0.015625,-0.0078125,0.015625,-0.015625,-0.0078125,0.03125,-0.0078125,-0.0,-0.046875,-0.03125,0.0078125,-0.0546875,-0.0234375,-0.0546875,-0.03125,0.0390625,-0.0078125,0.0546875,-0.0546875,0.0,0.0,0.0078125,0.015625,-0.0078125,0.0078125,0.0,0.0078125,-0.0078125,-0.0625,-0.0,-0.0078125,-0.09375,0.03125,0.0234375,0.015625,-0.0390625,-0.078125,0.0703125,0.0703125,0.046875,0.0234375,-0.015625,0.078125,-0.0390625,-0.03125,-0.0390625,0.0625,0.0625,-0.0546875,-0.0546875,-0.015625,0.0078125,-0.03125,-0.0390625,-0.046875,-0.03125,0.0390625,0.03125,-0.0390625,0.0078125,0.0625,-0.015625,-0.015625,-0.015625,-0.0234375,0.0078125,-0.0234375,-0.0,-0.0625,0.0390625,-0.0234375,-0.03125,-0.0390625,-0.0078125,-0.0546875,0.0390625,-0.0234375,0.0390625,-0.0078125,0.03125,0.0234375,-0.0,0.03125,0.0390625,-0.0078125,-0.0078125,0.0078125,0.0390625,-0.0234375,-0.015625,0.0,0.03125,0.0078125,-0.0234375,-0.03125,-0.0546875,-0.0234375,0.0234375,-0.0078125,0.0078125,-0.03125,-0.09375,-0.0,-0.0234375,-0.015625,0.0234375,0.0625,-0.0234375,-0.0625,0.015625,-0.0,0.078125,0.0078125,-0.0,-0.046875,0.015625,-0.0859375,-0.03125,-0.0,-0.0078125,-0.015625,-0.0078125,-0.0078125,-0.03125,0.0,0.0078125,0.0,-0.0078125,-0.0546875,-0.03125,0.0390625,0.046875,-0.03125,0.015625,-0.03125,-0.015625,-0.0234375,0.0234375,0.0234375,0.0,0.0078125,0.015625,-0.015625,-0.0,0.0078125,0.03125,-0.0,0.0859375,-0.0390625,-0.0234375,0.0625,-0.0234375,-0.015625,-0.0390625,-0.0,-0.0390625,0.046875,-0.078125,0.0078125,0.0078125,0.03125,0.0,-0.0234375,0.0234375,0.0,0.015625,-0.0390625,-0.0546875,-0.015625,-0.0390625,-0.0234375,-0.03125,0.0078125,0.0234375,-0.0390625,0.0390625,0.0625,0.0390625,-0.0390625,-0.015625,-0.0078125,0.046875,0.0234375,-0.015625,0.0859375,-0.046875,-0.0078125,-0.03125,0.015625,0.0,0.03125,-0.0625,0.015625,0.0625,0.015625,-0.0234375,0.03125,-0.0234375,-0.015625,0.0703125,-0.0,-0.0234375,0.09375,-0.046875,-0.0078125,-0.03125,-0.0234375,0.015625,-0.0390625,0.0078125,-0.0,-0.03125,-0.0625,-0.046875,-0.03125,-0.0078125,-0.0078125,-0.0859375,-0.03125,-0.0703125,-0.0234375,-0.0,-0.015625,0.0859375,0.03125,0.0078125,-0.0390625,0.078125,-0.0390625,0.0078125,-0.0078125,0.0625,-0.0234375,-0.0234375,-0.015625,-0.0390625,0.046875,-0.03125,0.03125,-0.0625,-0.0390625,-0.015625,-0.0390625,-0.015625,-0.0390625,0.0078125,0.0078125,-0.0,-0.0234375,0.0625,-0.015625,-0.0078125,0.046875,-0.0,0.0078125,-0.0,0.0625,-0.078125,0.0625,-0.015625,-0.0234375,-0.03125,0.0,0.0234375,0.0078125,-0.03125,0.0390625,0.0390625,-0.0625,0.0390625,0.0234375,-0.0078125,-0.0078125,-0.0078125,-0.0078125,-0.015625,-0.0078125,0.0,0.015625,-0.0078125,-0.03125,-0.0234375,0.0625,-0.0234375,-0.0703125,0.0078125,-0.0078125,0.0,0.0078125,-0.0234375,-0.015625,0.0078125,-0.0,-0.015625,0.046875,0.0234375,-0.0078125,0.0078125,0.109375,0.1015625,-0.0546875,-0.0234375,-0.0625,-0.015625,-0.0234375,-0.09375,0.015625,0.0078125,-0.0078125,-0.0078125,0.0,0.0078125,0.0078125,0.0,0.0078125,-0.015625,0.0390625,-0.0234375,0.0546875,0.0234375,-0.0234375,0.0234375,-0.0234375,0.015625,0.0,-0.0,0.078125,-0.015625,-0.0234375,-0.0625,-0.0625,-0.0078125,-0.015625,0.015625,0.09375,0.1171875,-0.03125,-0.109375,-0.0078125,-0.0078125,-0.0234375,-0.03125,0.015625,-0.0546875,-0.03125,0.0,-0.0234375,-0.0234375,-0.015625,0.0390625,0.0390625,-0.015625,-0.0234375,-0.03125,0.0,-0.0546875,-0.03125,-0.0078125,-0.0234375,-0.015625,-0.03125,0.015625,-0.0078125,-0.03125,0.015625,0.0,0.0234375,-0.0234375,0.0078125,0.015625,0.0546875,-0.0,-0.0546875,0.015625,0.03125,-0.0078125,-0.0,-0.0,0.0234375,0.03125,0.0234375,-0.0078125,-0.046875,0.0,0.0078125,0.0234375,0.0078125,0.0234375,-0.015625,0.03125,-0.046875,-0.0,-0.0703125,-0.0078125,-0.0234375,0.0234375,-0.0078125,-0.03125,0.046875,-0.015625,-0.0078125,0.015625,-0.0078125,-0.0078125,0.015625,-0.03125,-0.015625,-0.0,0.0,0.0,0.0078125,0.0078125,-0.0,0.015625,0.015625,0.0078125,-0.03125,0.0078125,0.0234375,-0.0,-0.015625,-0.015625,-0.0,-0.0,0.0078125,0.046875,0.0546875,-0.015625,-0.0078125,-0.0546875,-0.0234375,-0.015625,-0.03125,-0.015625,0.0625,-0.0234375,-0.03125,-0.046875,0.015625,0.015625,0.03125,-0.015625,0.046875,0.078125,0.0,-0.015625,-0.0625,-0.0625,0.0078125,-0.0078125,0.015625,-0.015625,-0.0859375,-0.1015625,0.015625,-0.015625,-0.03125,-0.0234375,0.0546875,-0.015625,0.0,-0.0546875,-0.03125,-0.015625,-0.015625,-0.0,-0.0390625,-0.03125,0.0078125,0.0625,0.0078125,-0.0390625,0.015625,-0.1015625,-0.0078125,0.0546875,0.0078125,0.0078125,-0.0234375,0.0078125,-0.015625,0.0703125,-0.046875,-0.0625,-0.03125,-0.046875,-0.015625,0.0859375,0.046875,-0.0390625,0.03125,-0.078125,-0.015625,-0.046875,-0.046875,0.0234375,0.0078125,0.0546875,-0.0078125,-0.0234375,0.03125,0.0,-0.0546875,0.0078125,0.0703125,0.140625,0.0078125,-0.015625,0.0078125,0.046875,0.0,-0.0390625,-0.03125,0.0234375,0.046875,-0.0859375,0.0546875,-0.046875,-0.0078125,-0.0625,0.015625,0.03125,-0.015625,-0.03125,-0.046875,-0.0078125,-0.015625,0.09375,-0.0234375,-0.015625,0.015625,-0.046875,-0.0234375,-0.015625,-0.015625,-0.015625,-0.0078125,-0.0078125,0.0234375,-0.0234375,-0.0390625,0.0078125,-0.03125,-0.0546875,-0.03125,0.0546875,-0.046875,-0.0390625,0.0,-0.0,0.0,-0.0078125,0.0078125,-0.0234375,0.015625,0.03125,-0.0078125,-0.0078125,-0.078125,0.0078125,-0.0,-0.0078125,-0.0078125,0.0078125,0.0078125,-0.0,-0.0078125,0.015625,-0.0078125,-0.0546875,-0.0,-0.0234375,-0.0390625,0.0390625,-0.015625,-0.0546875,0.015625,0.0078125,0.0078125,0.0,0.0078125,-0.0078125,0.0078125,-0.015625,-0.0390625,-0.0390625,0.0,0.0,0.03125,-0.015625,-0.0078125,0.03125,-0.015625,0.0234375,0.0078125,0.0078125,0.0,-0.015625,0.015625,-0.0078125,0.0078125,0.0,0.015625,-0.0078125,0.0078125,-0.015625,-0.0,0.0,-0.0078125,-0.0234375,-0.0234375,0.0625,-0.015625,-0.0234375,0.015625,0.046875,-0.0234375,-0.0390625,0.0390625,0.0,0.0234375,-0.0859375,-0.0234375,0.0234375,-0.0234375,-0.015625,-0.0546875,-0.03125,-0.0234375,-0.03125,0.015625,-0.0078125,-0.0390625,-0.015625,-0.0,-0.0390625,0.0703125,-0.015625,-0.0,-0.0234375,0.015625,0.015625,0.03125,-0.0078125,-0.0390625,-0.0390625,-0.0,0.046875,0.0,0.015625,-0.0390625,0.015625,-0.015625,0.0390625,0.015625,-0.0078125,0.0078125,-0.046875,0.0078125,0.0,0.0390625,-0.0,-0.0078125,-0.015625,-0.0,0.015625,-0.0,-0.0078125,0.0,0.0,-0.015625,-0.015625,0.015625,-0.0234375,0.0078125,0.015625,-0.0078125,-0.046875,-0.03125,-0.0234375,-0.0234375,-0.0078125,0.0078125,0.0625,0.03125,0.0,0.0,-0.0234375,-0.015625,0.0078125,-0.0390625,-0.0078125,0.0234375,0.0390625,0.0078125,0.0078125,0.0,-0.0078125,0.015625,0.0078125,0.0,-0.0078125,0.0234375,0.0,-0.03125,-0.0,-0.015625,-0.0078125,0.0,-0.0,-0.0,0.03125,0.0078125,0.0,-0.0078125,0.0,-0.0078125,-0.046875,-0.0078125,0.0703125,0.0078125,-0.015625,-0.0390625,-0.0625,0.015625,-0.0390625,0.046875,-0.0078125,-0.0,0.015625,-0.0078125,0.015625,-0.0,-0.0078125,-0.0390625,-0.109375,-0.0234375,0.03125,0.046875,-0.0078125,0.0390625,0.0234375,-0.015625,-0.0,-0.078125,-0.03125,0.015625,0.046875,0.0078125,0.0078125,-0.0,0.0,0.015625,0.015625,-0.0234375,-0.0546875,-0.0,-0.015625,-0.015625,-0.046875,-0.015625,0.015625,0.0625,0.0,-0.09375,-0.015625,-0.0078125,-0.03125,-0.0390625,-0.0078125,-0.0078125,0.03125,0.0078125,-0.015625,0.046875,-0.0078125,0.0390625,0.0234375,-0.0078125,-0.0234375,-0.046875,0.0,-0.0703125,-0.015625,-0.0,-0.0703125,0.078125,0.0,-0.0078125,-0.046875,-0.0234375,0.03125,-0.0234375,-0.015625,-0.0078125,-0.0546875,-0.03125,0.0390625,-0.09375,-0.015625,0.0,0.0390625,-0.015625,-0.0078125,0.015625,-0.0,0.015625,-0.0,-0.0078125,0.0625,0.0390625,-0.0078125,-0.046875,0.0234375,-0.015625,0.0234375,0.0078125,-0.0078125,-0.03125,-0.0625,-0.0,-0.0078125,0.046875,-0.015625,0.0625,0.0703125,-0.0234375,-0.015625,0.0234375,0.0078125,0.0546875,0.0390625,-0.015625,0.0234375,0.0,-0.015625,-0.0390625,-0.015625,-0.0234375,0.0234375,-0.0234375,-0.03125,0.0625,0.0234375,0.0625,0.0234375,-0.0078125,-0.0078125,-0.0,0.0,0.0078125,-0.0078125,-0.0078125,-0.0078125,-0.0078125,0.0,0.046875,0.03125,-0.0234375,0.015625,-0.015625,0.0,0.0234375,0.0390625,-0.015625,0.0078125,-0.0390625,-0.0546875,0.0234375,-0.1015625,0.0234375,-0.0625,0.046875,-0.03125,0.0703125,0.0703125,-0.015625,0.03125,-0.0390625,0.0234375,0.0703125,-0.0390625,-0.03125,-0.0,0.0078125,0.0,0.015625,-0.0078125,0.0078125,-0.0078125,-0.0078125,-0.0,-0.015625,0.046875,-0.03125,0.0,-0.0859375,-0.03125,-0.0078125,-0.0859375,-0.03125,0.0546875,-0.0,-0.0,-0.0234375,0.0390625,-0.0078125,0.0234375,0.0078125,-0.0234375,0.0234375,0.046875,-0.0234375,0.015625,-0.0,0.0234375,0.0078125,-0.046875,-0.0390625,-0.046875,0.0546875,0.015625,-0.015625,0.015625,0.0078125,-0.015625,-0.0234375,-0.0078125,0.0703125,0.03125,-0.0703125,-0.03125,0.0078125,-0.0234375,-0.0,0.0234375,-0.0234375,-0.015625,0.0,0.0390625,0.0390625,-0.015625,-0.0078125,-0.0,-0.03125,0.0,0.0234375,-0.0078125,-0.015625,-0.0,0.0078125,-0.0234375,0.0,-0.015625,-0.0,0.0,-0.015625,0.0625,-0.0390625,-0.0625,-0.0078125,-0.0390625,0.015625,-0.015625,0.0078125,0.046875,-0.03125,-0.0078125,0.0078125,-0.0390625,-0.015625,-0.03125,-0.0,0.0234375,0.0078125,0.015625,0.0625,-0.0078125,-0.015625,-0.015625,-0.0859375,-0.015625,0.015625,-0.0078125,-0.0078125,-0.015625,0.015625,0.0078125,0.0078125,-0.0,-0.015625,-0.0078125,-0.0703125,-0.0078125,-0.0625,-0.03125,-0.0234375,0.0078125,-0.015625,-0.0078125,-0.0078125,-0.0390625,0.0078125,-0.0546875,0.046875,-0.015625,-0.0546875,0.0546875,-0.0390625,0.0,0.0546875,0.0,0.0625,-0.0234375,0.0390625,-0.03125,-0.0546875,0.0078125,-0.03125,0.0078125,-0.0390625,-0.015625,-0.0234375,-0.0390625,-0.046875,-0.0078125,-0.015625,0.046875,-0.0546875,-0.0390625,-0.1015625,-0.0078125,-0.0,-0.0625,-0.0234375,-0.0234375,0.0,0.015625,-0.015625,0.015625,0.046875,-0.0234375,0.046875,0.046875,-0.015625,-0.0546875,-0.078125,0.0546875,0.0546875,-0.015625,0.0,0.03125,0.0,-0.0390625,-0.0078125,-0.0546875,-0.0078125,-0.0078125,-0.0234375,-0.0234375,0.0625,-0.0625,-0.0,-0.03125,-0.015625,-0.0078125,-0.0390625,-0.015625,-0.03125,0.171875,-0.0234375,-0.0078125,-0.015625,0.0078125,-0.0,0.0390625,-0.0625,0.0859375,0.0234375,0.0234375,-0.03125,-0.0390625,-0.0625,0.1015625,-0.0703125,0.03125,-0.0546875,0.0,0.0234375,-0.03125,-0.0546875,-0.03125,-0.015625,0.0,-0.078125,-0.0390625,-0.0703125,-0.0703125,-0.015625,-0.0078125,0.0078125,-0.0390625,-0.046875,-0.0546875,-0.0078125,-0.0703125,0.0390625,-0.0234375,0.0,-0.0078125,-0.015625,0.046875,0.0859375,-0.0078125,-0.015625,-0.015625,0.0,-0.1171875,0.015625,-0.03125,-0.0625,-0.0546875,-0.0078125,-0.0,0.046875,-0.015625,0.0390625,0.0078125,0.078125,-0.03125,-0.015625,-0.0078125,0.03125,-0.0,0.0703125,-0.0078125,-0.0078125,-0.0078125,0.015625,0.0,0.0078125,-0.0078125,0.015625,-0.0078125,0.015625,-0.0078125,-0.1328125,-0.03125,-0.015625,-0.1015625,0.0390625,-0.0078125,0.0234375,0.0078125,0.0234375,-0.015625,-0.015625,0.046875,-0.0859375,0.0546875,0.0234375,0.0,-0.0234375,0.0078125,0.03125,-0.0078125,-0.078125,-0.0,-0.0390625,-0.0390625,-0.0390625,0.0,-0.015625,-0.0078125,-0.0,0.015625,0.0,0.0,-0.0078125,-0.0078125,-0.03125,-0.0234375,-0.046875,-0.046875,0.03125,-0.0234375,-0.03125,-0.03125,-0.0078125,0.078125,0.0390625,-0.0234375,0.0390625,-0.0390625,-0.0703125,-0.015625,0.0390625,0.0625,-0.0234375,-0.0703125,-0.0390625,0.0,-0.0234375,0.03125,-0.0234375,-0.03125,0.046875,-0.0,0.0234375,-0.015625,-0.0078125,-0.0234375,0.0234375,0.0234375,0.0,0.0234375,-0.0078125,-0.015625,0.0703125,0.0078125,-0.03125,-0.03125,-0.015625,0.0390625,0.03125,-0.0,0.0,0.0,-0.015625,-0.015625,-0.046875,-0.03125,0.015625,0.0390625,-0.015625,-0.0390625,-0.0078125,0.0,-0.0078125,-0.03125,-0.015625,0.0390625,0.0234375,-0.0078125,-0.078125,-0.0078125,0.0234375,-0.0078125,0.0234375,-0.0,-0.03125,-0.0703125,-0.0,0.1015625,0.1015625,0.0,-0.0078125,-0.0703125,-0.0,0.0703125,-0.0234375,-0.015625,-0.0234375,-0.0078125,0.0234375,-0.0078125,0.125,0.0078125,-0.015625,-0.046875,0.0,-0.015625,-0.0078125,0.0,0.0078125,0.015625,0.0,0.0078125,-0.015625,-0.0078125,0.0,-0.0234375,-0.015625,0.015625,0.0,-0.015625,-0.0234375,0.046875,0.03125,0.0546875,0.015625,0.015625,0.03125,0.0,-0.0234375,0.1015625,-0.015625,0.0078125,0.015625,0.109375,0.015625,-0.0703125,-0.046875,-0.0,-0.0,0.0703125,-0.0078125,0.0234375,0.1015625,-0.0234375,0.0390625,-0.0390625,-0.0234375,0.015625,-0.046875,-0.0078125,0.015625,0.015625,-0.0078125,-0.0078125,0.03125,-0.0390625,-0.03125,0.09375,0.0234375,-0.0234375,-0.0234375,-0.0546875,-0.0,0.0078125,-0.0078125,0.015625,-0.0234375,0.015625,0.0546875,0.0,0.015625,-0.0078125,-0.0625,0.0390625,0.0234375,-0.0234375,-0.03125,-0.0390625,0.046875,-0.015625,-0.0234375,0.09375,-0.015625,0.03125,0.0234375,0.0234375,0.0234375,0.015625,-0.0,-0.046875,-0.0078125,0.0,-0.0703125,-0.0703125,0.0234375,-0.0234375,0.0390625,-0.0078125,0.0390625,0.03125,-0.015625,0.015625,-0.0234375,-0.046875,-0.0234375,0.03125,-0.0390625,-0.078125,-0.015625,0.0,-0.0078125,-0.03125,-0.0078125,-0.03125,0.0625,0.015625,-0.015625,-0.109375,0.0234375,-0.015625,0.0234375,0.0,-0.0078125,-0.09375,-0.015625,-0.0546875,-0.0625,0.015625,0.03125,-0.0625,0.0625,-0.0859375,0.0390625,-0.046875,-0.0078125,-0.015625,-0.0078125,-0.015625,-0.0234375,0.03125,0.125,-0.0703125,-0.0078125,-0.0625,-0.015625,-0.0234375,-0.0,-0.046875,-0.0234375,-0.015625,0.0390625,-0.0234375,0.0234375,0.015625,0.015625,-0.0234375,-0.015625,0.0078125,-0.0078125,0.0078125,0.0,0.0,0.0078125,-0.0,0.015625,0.015625,-0.015625,-0.0625,0.03125,-0.078125,-0.0390625,0.0703125,0.0078125,-0.03125,-0.0234375,0.03125,-0.03125,0.0234375,0.0078125,-0.046875,0.0703125,-0.015625,-0.0078125,0.0078125,-0.0,0.0234375,0.0,-0.046875,0.03125,0.078125,-0.0234375,-0.0,-0.046875,-0.0,0.0,-0.015625,0.0078125,-0.0,0.0078125,-0.0078125,-0.0078125,-0.0078125,0.0625,-0.0546875,0.09375,-0.0625,-0.0859375,0.0234375,-0.03125,-0.046875,-0.0078125,0.0078125,0.0390625,0.0546875,-0.015625,0.0078125,0.03125,-0.0078125,-0.0234375,0.0078125,-0.0078125,0.0859375,0.015625,-0.0390625,0.0234375,-0.109375,-0.03125,-0.046875,-0.0234375,0.03125,-0.03125,-0.0,-0.0078125,0.0234375,-0.0078125,-0.015625,-0.0390625,-0.0,0.0625,-0.03125,-0.0703125,-0.0078125,0.0078125,0.015625,0.0078125,-0.0234375,0.0078125,-0.0234375,0.015625,0.03125,-0.046875,-0.0234375,-0.0234375,0.0078125,-0.0,-0.0,0.015625,-0.0,-0.015625,0.0078125,-0.015625,-0.0234375,0.0,0.0,-0.0078125,-0.015625,0.046875,-0.0625,-0.0078125,-0.015625,-0.046875,0.0,0.0234375,0.0234375,0.03125,-0.0078125,-0.0625,0.0078125,0.0234375,0.03125,-0.0,-0.03125,-0.015625,-0.03125,0.0859375,-0.015625,-0.078125,0.03125,-0.03125,-0.0234375,-0.0234375,-0.015625,-0.015625,0.015625,-0.015625,-0.0,0.0078125,0.0234375,-0.0078125,-0.0,-0.0,0.0,-0.0078125,0.0078125,-0.0625,-0.0390625,0.0546875,0.015625,-0.0234375,0.0234375,0.0390625,-0.0703125,-0.0,0.03125,-0.03125,0.0078125,-0.0078125,-0.015625,0.0,0.0078125,0.0390625,0.0625,-0.0234375,0.0390625,-0.0546875,-0.0234375,0.0078125,-0.0078125,-0.015625,0.03125,0.0,-0.0078125,-0.046875,-0.0,-0.0078125,0.0078125,0.03125,-0.0703125,-0.046875,-0.0,-0.0703125,0.0390625,0.046875,0.0234375,0.015625,-0.015625,0.015625,0.0703125,0.046875,0.0234375,-0.046875,-0.0078125,-0.0234375,-0.0078125,-0.0078125,-0.0390625,0.0078125,-0.0625,0.0234375,-0.03125,-0.0234375,0.015625,-0.015625,0.0078125,-0.0546875,0.0234375,-0.0234375,-0.0234375,-0.0078125,0.0390625,-0.015625,-0.0,0.03125,-0.03125,0.046875,-0.0546875,-0.0078125,-0.0,-0.0546875,0.0234375,0.0078125,0.0,0.0,-0.015625,-0.015625,-0.0078125,0.078125,-0.0234375,0.0078125,-0.0078125,-0.0390625,0.078125,0.0546875,0.0078125,0.015625,-0.0859375,-0.078125,-0.0078125,-0.0390625,-0.0,0.0078125,-0.078125,-0.03125,0.03125,0.09375,0.03125,-0.0234375,0.0234375,0.0,0.015625,-0.0859375,-0.0390625,-0.0390625,-0.0390625,0.03125,0.0078125,-0.0078125,-0.0234375,-0.0,0.0234375,0.0234375,-0.03125,-0.0078125,0.0625,0.015625,-0.0234375,0.0,0.0859375,-0.0234375,0.0390625,0.0078125,-0.015625,0.0078125,0.0078125,-0.015625,-0.0,-0.0390625,-0.0546875,-0.03125,-0.0078125,-0.046875,0.09375,-0.0234375,-0.0078125,0.0078125,-0.0078125,-0.0,-0.0078125,0.0,0.0078125,0.0078125,0.015625,-0.0078125,0.0234375,-0.0625,0.03125,0.03125,-0.0078125,0.046875,-0.015625,-0.015625,-0.0,-0.0,-0.046875,-0.03125,0.0078125,0.0078125,0.078125,0.046875,-0.0078125,-0.0,-0.0,-0.0078125,-0.015625,-0.0390625,0.0,-0.0234375,-0.0234375,0.015625,0.0625,-0.0234375,0.0,0.0078125,-0.015625,0.015625,-0.015625,0.0,0.0,-0.0078125,-0.0078125,-0.0390625,0.03125,-0.03125,-0.0234375,-0.0703125,-0.0390625,-0.0234375,-0.0078125,0.03125,-0.0390625,0.015625,-0.0625,-0.015625,-0.0390625,0.0859375,-0.03125,-0.0703125,-0.046875,-0.0078125,-0.0625,-0.0078125,-0.015625,0.0,-0.0390625,-0.0625,-0.015625,-0.0859375,-0.0,0.015625,-0.0078125,-0.0390625,-0.0546875,-0.0703125,-0.0234375,0.0078125,-0.0390625,-0.0234375,-0.0859375,-0.0546875,-0.046875,-0.015625,-0.03125,0.0078125,0.015625,0.0390625,0.0078125,-0.0078125,-0.015625,0.046875,-0.0,-0.03125,0.0078125,-0.0546875,0.03125,0.0234375,0.078125,0.0078125,-0.0,-0.0234375,-0.0234375,-0.0078125,0.0078125,0.0078125,-0.0,0.0234375,-0.0234375,0.015625,-0.0390625,-0.0390625,-0.0234375,0.015625,-0.0078125,-0.03125,-0.046875,-0.03125,-0.0234375,-0.078125,0.078125,-0.0078125,-0.0078125,-0.03125,-0.0078125,-0.0234375,-0.0859375,-0.0546875,-0.0234375,0.0234375,-0.0,0.03125,-0.0234375,0.0078125,0.0,0.015625,0.015625,-0.0,0.0,-0.015625,0.0,0.015625,-0.0078125,0.0546875,-0.03125,0.015625,0.0390625,-0.0078125,-0.0234375,0.0078125,0.0078125,-0.0,0.03125,-0.0,-0.015625,-0.015625,-0.0390625,0.0,0.0546875,0.0078125,-0.0078125,-0.03125,0.03125,0.0390625,0.0390625,0.015625,0.015625,-0.03125,-0.0234375,0.0546875,-0.0546875,0.0390625,-0.046875,-0.0625,0.0234375,-0.0234375,-0.0546875,0.015625,-0.0078125,0.1015625,-0.0078125,0.0078125,-0.0078125,-0.046875,0.0234375,0.0625,-0.0859375,-0.0,0.09375,0.0390625,-0.03125,0.0234375,-0.0625,-0.0234375,0.0078125,-0.0234375,-0.0,0.09375,-0.0234375,0.0,-0.0078125,0.0078125,0.0,0.0234375,0.0234375,0.0,-0.0234375,0.0078125,0.0,-0.0078125,-0.0078125,0.0234375,-0.0078125,0.03125,0.0390625,0.03125,-0.0390625,0.0390625,-0.0078125,-0.015625,-0.0078125,-0.015625,0.0234375,-0.0234375,0.1015625,-0.0234375,-0.0078125,0.046875,0.03125,0.0390625,-0.0,0.0234375,-0.03125,0.0546875,-0.0390625,-0.078125,-0.0625,0.015625,-0.03125,0.0078125,0.03125,-0.0234375,-0.0078125,0.0390625,-0.0234375,-0.046875,0.015625,0.0234375,-0.0078125,0.0546875,-0.0390625,0.15625,-0.0390625,-0.015625,-0.0234375,-0.0546875,-0.0234375,0.1015625,0.0546875,-0.03125,0.015625,-0.0234375,-0.0078125,-0.03125,-0.015625,-0.0078125,-0.015625,0.0234375,-0.0234375,0.015625,-0.0546875,-0.03125,0.015625,0.046875,-0.0390625,-0.0,-0.015625,-0.03125,-0.046875,-0.03125,-0.0078125,-0.015625,0.015625,0.0625,0.0546875,-0.03125,0.0078125,-0.0078125,-0.015625,-0.0078125,-0.0078125,-0.0078125,-0.0,-0.0,-0.0078125,-0.046875,0.0234375,0.046875,-0.0625,-0.0546875,0.0078125,0.03125,0.09375,-0.09375,0.015625,-0.0546875,0.0546875,0.015625,-0.0078125,-0.0234375,0.0625,0.0859375,-0.0390625,0.1015625,0.0078125,0.0390625,-0.0703125,-0.0078125,-0.0390625,-0.046875,0.0078125,-0.0234375,-0.0078125,-0.0078125,0.015625,0.0,-0.0078125,0.0,-0.0078125,0.0,-0.0078125,0.0625,-0.046875,-0.0078125,0.140625,-0.0,-0.0625,0.078125,0.0078125,0.015625,0.0703125,0.03125,0.0703125,0.0078125,0.0078125,-0.0390625,0.0,-0.015625,-0.0078125,0.0078125,-0.0625,-0.0,-0.0234375,-0.03125,-0.0625,0.046875,0.0078125,-0.03125,0.0,0.015625,-0.015625,0.0625,0.046875,0.0078125,-0.0390625,-0.03125,-0.0078125,0.0234375,-0.0234375,-0.015625,-0.0078125,-0.03125,0.0078125,-0.015625,-0.078125,-0.015625,0.0234375,-0.0234375,-0.03125,-0.0625,0.0,0.0390625,0.0234375,-0.015625,0.0078125,0.03125,0.0546875,0.03125,-0.0234375,0.015625,0.015625,-0.015625,-0.015625,0.015625,0.0,-0.015625,0.0234375,-0.0546875,-0.015625,0.0078125,-0.0234375,0.015625,-0.015625,0.046875,0.015625,-0.015625,0.0234375,-0.0546875,-0.03125,-0.0078125,-0.0546875,-0.0546875,0.0703125,0.125,-0.078125,-0.015625,-0.09375,-0.015625,-0.0625,-0.0,-0.078125,-0.0078125,-0.015625,0.0078125,0.0078125,-0.015625,-0.0078125,-0.015625,-0.0,-0.0,0.015625,-0.0,-0.015625,-0.0078125,-0.0546875,0.015625,0.0625,-0.0234375,-0.03125,-0.0078125,-0.0234375,-0.0078125,-0.0078125,0.0234375,0.0390625,0.0,0.0390625,-0.03125,-0.0078125,0.0390625,0.0390625,0.046875,-0.03125,-0.0390625,-0.0234375,0.015625,-0.0234375,0.0,-0.015625,0.0234375,0.0,-0.0234375,0.015625,-0.03125,-0.03125,0.015625,-0.03125,0.0625,0.0078125,0.03125,-0.0546875,-0.0234375,-0.015625,-0.0546875,0.0390625,-0.0,-0.0078125,0.0390625,-0.0390625,-0.046875,0.0,0.0625,0.09375,0.0,0.0546875,-0.0390625,0.03125,-0.0546875,-0.0625,0.078125,0.0,0.0078125,-0.0078125,-0.0,-0.0078125,-0.046875,0.0,-0.046875,0.0,0.0390625,-0.0390625,-0.0234375,-0.0390625,-0.0546875,-0.0,-0.0390625,0.0625,0.015625,-0.03125,-0.0,0.0703125,-0.0078125,0.0859375,0.03125,-0.0234375,-0.0234375,-0.0703125,0.046875,0.0546875,0.03125,0.0234375,-0.0078125,-0.0625,0.0078125,-0.09375,0.015625,0.0078125,-0.0234375,0.0078125,0.1484375,-0.015625,-0.0078125,-0.0234375,-0.0703125,-0.046875,-0.0390625,-0.046875,-0.078125,-0.03125,0.0,-0.0,-0.0078125,-0.03125,-0.015625,-0.046875,0.0,-0.0,0.046875,0.1328125,0.0546875,-0.109375,0.0234375,-0.015625,-0.0,-0.015625,-0.03125,-0.015625,-0.0546875,-0.0234375,-0.046875,-0.0234375,-0.0234375,0.0,-0.015625,0.0,0.0078125,0.0234375,0.0078125,0.0078125,-0.0703125,0.0,-0.015625,0.0078125,0.0859375,-0.0,0.0,-0.0078125,-0.015625,0.0078125,0.0078125,-0.0078125,0.0,-0.0,0.015625,-0.0234375,-0.015625,-0.0078125,0.0234375,0.046875,0.0,-0.0078125,-0.0234375,-0.0078125,0.0234375,0.0,0.0,0.0078125,0.0,-0.0078125,-0.0234375,-0.0234375,-0.0234375,-0.0625,-0.0078125,-0.0390625,0.046875,0.0546875,-0.0234375,-0.0390625,-0.046875,0.0078125,-0.0078125,-0.0078125,0.0,-0.0078125,-0.0078125,-0.0078125,0.0078125,0.0078125,-0.03125,0.0234375,0.03125,-0.0390625,-0.03125,-0.078125,0.0,-0.0390625,0.015625,-0.015625,0.078125,-0.046875,-0.0234375,0.0234375,0.015625,-0.0234375,0.046875,-0.015625,0.015625,0.078125,0.0,-0.0546875,-0.0078125,0.0546875,-0.0390625,-0.046875,-0.078125,0.0390625,0.03125,0.0078125,0.03125,-0.03125,0.0,-0.015625,-0.03125,-0.0234375,-0.015625,0.0078125,0.046875,-0.03125,0.0,-0.015625,-0.0234375,-0.0234375,-0.0234375,-0.03125,-0.0234375,-0.0234375,-0.015625,0.03125,-0.0078125,-0.0078125,-0.015625,-0.015625,-0.0234375,-0.015625,-0.015625,-0.015625,-0.03125,0.0078125,0.0078125,0.0078125,-0.0078125,-0.0234375,0.0,0.015625,-0.0,0.015625,0.03125,-0.015625,0.015625,-0.0234375,0.0,-0.03125,0.0390625,-0.0078125,-0.0078125,-0.0390625,-0.0078125,-0.0234375,-0.0078125,-0.015625,-0.015625,-0.0078125,-0.015625,-0.0078125,-0.0078125,-0.03125,0.0,0.0390625,-0.0078125,0.015625,0.0,-0.0078125,-0.0,0.0078125,-0.0078125,0.0234375,0.0078125,-0.03125,-0.046875,0.0078125,-0.0078125,0.015625,0.015625,-0.0,-0.0078125,0.015625,0.015625,0.0,-0.0234375,-0.0078125,0.0234375,0.0078125,-0.015625,-0.015625,-0.0234375,0.03125,0.0703125,0.0234375,-0.03125,0.0078125,0.0859375,-0.015625,-0.0390625,-0.078125,-0.0546875,-0.015625,-0.0546875,0.0,0.0546875,0.0390625,-0.015625,-0.0234375,0.0546875,-0.015625,0.0078125,0.0078125,-0.0078125,-0.0859375,0.0546875,0.0078125,-0.03125,-0.0390625,0.015625,-0.0,-0.03125,-0.0234375,0.0390625,0.015625,-0.0234375,-0.0234375,-0.015625,0.015625,-0.0234375,-0.015625,0.0078125,-0.0078125,0.0546875,-0.015625,0.0390625,-0.0625,-0.0234375,0.0078125,0.0,-0.015625,0.046875,0.0546875,-0.0078125,-0.0546875,-0.015625,-0.046875,0.015625,-0.046875,-0.0234375,0.0703125,-0.03125,-0.0078125,-0.03125,-0.015625,-0.0,-0.0078125,-0.015625,-0.078125,-0.09375,-0.0546875,-0.0078125,-0.0078125,0.046875,0.0078125,-0.0703125,-0.0703125,-0.015625,0.0390625,0.0390625,-0.0078125,-0.0625,-0.046875,-0.0078125,-0.0078125,-0.0390625,-0.0,0.046875,-0.046875,-0.0078125,-0.015625,-0.0078125,-0.0546875,-0.03125,-0.015625,-0.0234375,-0.03125,-0.09375,-0.0078125,-0.0390625,0.0390625,-0.0078125,-0.0703125,-0.0703125,-0.0390625,0.03125,-0.0078125,-0.0234375,0.015625,0.15625,-0.0234375,-0.0,-0.03125,-0.0234375,0.015625,-0.0234375,-0.0234375,0.0390625,-0.0390625,0.0234375,-0.03125,-0.0390625,0.0078125,-0.0,-0.015625,0.0390625,0.09375,-0.0078125,0.0078125,-0.015625,-0.0,-0.0,-0.0,-0.0234375,0.0,-0.0078125,0.0,-0.015625,0.0625,-0.046875,-0.0546875,-0.1015625,-0.078125,-0.0078125,0.1015625,0.0234375,0.0078125,0.078125,-0.0234375,0.03125,-0.03125,-0.015625,0.0390625,-0.015625,-0.03125,0.03125,-0.0078125,0.03125,-0.0703125,-0.0234375,-0.046875,-0.078125,0.0078125,0.03125,-0.0,-0.015625,-0.0078125,-0.0078125,-0.0,0.0078125,0.0078125,0.0,0.0078125,0.0234375,0.0078125,0.0390625,0.03125,0.03125,-0.03125,-0.0625,0.0546875,0.0,0.0078125,0.1484375,-0.0625,-0.0078125,-0.09375,-0.078125,0.015625,0.0078125,-0.03125,0.015625,-0.0078125,0.0078125,0.0078125,-0.0078125,0.015625,0.015625,-0.0078125,0.0078125,0.0234375,-0.0,0.0078125,0.015625,0.0078125,0.0546875,0.0234375,-0.03125,0.0234375,-0.0,-0.0234375,0.0546875,0.0,0.015625,-0.015625,-0.0625,0.015625,-0.0390625,-0.015625,0.015625,0.0234375,-0.0,0.0078125,-0.0078125,-0.0234375,-0.03125,-0.0625,-0.0,0.0703125,0.0078125,-0.0390625,-0.0234375,-0.0390625,-0.03125,-0.0078125,-0.015625,0.0078125,-0.015625,-0.015625,0.03125,-0.03125,-0.0078125,-0.046875,-0.0390625,-0.015625,-0.015625,-0.0234375,-0.0,0.0078125,0.109375,0.0390625,-0.0078125,-0.0390625,0.0,0.0546875,0.046875,0.0078125,-0.0078125,-0.0234375,-0.015625,0.0078125,-0.0,0.0078125,0.0078125,-0.0,0.0078125,0.0,-0.0234375,-0.0078125,0.0078125,0.0078125,0.015625,0.0,0.125,-0.015625,-0.03125,0.046875,-0.0390625,-0.0078125,0.03125,0.0,-0.0390625,0.0625,-0.015625,-0.0234375,-0.0234375,0.0,-0.03125,-0.0390625,-0.0078125,-0.046875,-0.125,0.0234375,-0.0234375,0.03125,-0.03125,0.0390625,0.0703125,0.0546875,0.0234375,-0.03125,0.0703125,-0.03125,-0.0859375,-0.0859375,-0.0390625,-0.09375,-0.015625,-0.046875,-0.015625,-0.078125,-0.046875,-0.046875,-0.0546875,-0.0078125,0.0,-0.0234375,0.0,-0.0078125,-0.0234375,-0.0703125,-0.0234375,0.0390625,-0.015625,-0.03125,0.015625,-0.0078125,0.03125,-0.046875,-0.03125,-0.0859375,-0.0,0.03125,-0.046875,-0.03125,0.0390625,-0.0390625,0.03125,-0.0390625,0.03125,-0.03125,-0.0,-0.0078125,-0.0703125,-0.0078125,-0.0703125,-0.015625,-0.0546875,-0.0078125,-0.078125,0.0078125,-0.0703125,-0.0859375,0.046875,-0.015625,0.0078125,-0.0234375,-0.046875,-0.0234375,0.0234375,0.015625,0.0078125,-0.046875,0.1015625,-0.03125,0.0078125,-0.0234375,-0.0078125,-0.015625,-0.078125,-0.0234375,0.0078125,-0.078125,0.015625,0.0546875,0.0546875,-0.0,-0.078125,-0.078125,-0.0625,-0.046875,0.0546875,-0.03125,-0.015625,-0.03125,0.0078125,-0.0546875,-0.109375,0.0078125,0.0546875,0.0234375,0.046875,-0.03125,-0.0859375,-0.03125,-0.0234375,-0.015625,-0.0390625,-0.03125,0.0859375,-0.0390625,-0.0234375,-0.0859375,0.0,-0.015625,0.0234375,0.0,-0.015625,-0.078125,0.046875,0.0078125,-0.015625,0.0625,0.046875,0.015625,-0.0234375,0.015625,0.0078125,0.0,0.0,-0.0078125,0.015625,-0.0078125,-0.0234375,-0.0234375,-0.015625,-0.03125,-0.0546875,-0.0078125,0.03125,-0.1015625,0.0625,0.0234375,-0.0234375,-0.0078125,-0.03125,-0.0390625,0.1015625,-0.0546875,-0.0546875,0.0234375,-0.0234375,-0.0546875,0.0078125,-0.0,-0.015625,-0.0859375,-0.0625,0.0859375,-0.0390625,-0.0625,-0.046875,0.0,-0.015625,0.0078125,-0.0078125,0.0078125,-0.015625,-0.015625,-0.0078125,-0.0,0.0,0.0234375,0.015625,-0.015625,-0.0,-0.046875,-0.03125,0.0078125,-0.046875,0.015625,-0.0546875,0.078125,-0.015625,-0.046875,0.09375,-0.0234375,-0.0859375,0.03125,-0.0078125,-0.0859375,0.015625,-0.03125,-0.015625,0.03125,-0.046875,0.0078125,-0.03125,0.015625,-0.0078125,0.046875,-0.015625,0.015625,-0.03125,0.03125,0.03125,0.0390625,0.078125,0.0703125,0.078125,-0.0234375,-0.03125,0.0,0.0,0.015625,0.0,-0.0078125,-0.0,-0.0,0.0078125,0.0234375,0.09375,-0.0234375,-0.015625,0.0078125,-0.015625,-0.0234375,0.0078125,0.0078125,0.046875,0.0078125,-0.015625,0.0078125,0.0078125,0.0234375,0.015625,-0.015625,0.0078125,0.0078125,-0.0234375,-0.0234375,-0.0,0.03125,-0.0234375,-0.03125,0.125,0.078125,-0.046875,-0.03125,0.03125,-0.0078125,0.015625,0.0078125,0.0234375,0.0078125,-0.015625,-0.0078125,0.046875,-0.0078125,-0.0234375,-0.03125,-0.015625,-0.015625,-0.0078125,0.0078125,-0.03125,0.0078125,0.0078125,-0.0078125,0.0,0.0078125,-0.0546875,0.03125,-0.0078125,0.03125,0.0625,0.0,0.0625,-0.046875,0.078125,-0.0234375,-0.015625,-0.0234375,0.015625,-0.03125,0.0390625,0.0234375,0.03125,0.03125,0.015625,0.0234375,-0.0390625,-0.078125,0.0234375,-0.015625,-0.0078125,0.09375,0.0078125,-0.0390625,-0.03125,-0.125,0.0546875,-0.046875,0.046875,0.0546875,0.0234375,0.0,-0.0,-0.046875,-0.0625,-0.0234375,0.078125,-0.0,-0.0234375,0.015625,-0.0703125,-0.078125,-0.03125,0.0390625,0.015625,-0.0,0.046875,-0.0703125,0.0703125,0.0703125,0.140625,-0.0703125,-0.0703125,-0.0703125,-0.140625,0.0703125,-0.0234375,0.0390625,-0.0234375,-0.0546875,0.0234375,-0.0390625,-0.0,0.1015625,0.0390625,-0.03125,-0.03125,-0.078125,-0.0234375,-0.0078125,-0.0234375,0.125,-0.0703125,0.03125,-0.09375,-0.078125,0.0625,0.0390625,-0.0703125,-0.046875,0.0078125,0.0078125,0.015625,0.0234375,-0.046875,0.0625,0.0390625,0.1171875,-0.046875,-0.0546875,-0.0625,-0.015625,0.078125,0.0546875,0.1015625,-0.0078125,0.046875,-0.0390625,-0.0078125,0.0078125,0.0703125,0.0078125,0.078125,0.046875,0.0625,-0.0234375,0.015625,-0.0234375,0.0,-0.0625,-0.0390625,-0.015625,-0.03125,-0.0078125,-0.0546875,-0.0,0.0703125,-0.0390625,-0.015625,-0.046875,-0.0390625,0.0390625,0.0078125,0.015625,-0.03125,-0.0234375,-0.0390625,0.0546875,-0.0546875,-0.0234375,0.0078125,-0.046875,-0.0234375,-0.0,-0.046875,-0.0234375,0.078125,0.0234375,0.0234375,0.015625,-0.0078125,-0.015625,-0.0,0.0078125,-0.0078125,-0.0,-0.0078125,0.0,-0.0078125,0.15625,-0.0234375,-0.046875,-0.0625,-0.03125,0.0,-0.0078125,0.015625,0.0390625,-0.0078125,0.0078125,0.0,-0.046875,-0.046875,-0.0,-0.015625,0.03125,0.015625,-0.0,-0.03125,0.0,-0.0546875,-0.1015625,-0.0546875,0.0703125,-0.0390625,0.0078125,0.0,0.0,0.0,0.0078125,0.0,0.0078125,0.015625,0.0078125,-0.0234375,0.03125,0.0234375,-0.046875,-0.03125,-0.078125,-0.0546875,0.03125,-0.0078125,0.0,0.046875,0.0234375,0.03125,-0.0546875,-0.0546875,0.046875,0.0078125,0.0234375,-0.0390625,-0.0,-0.0390625,-0.0546875,0.0859375,0.109375,0.078125,-0.03125,0.0546875,-0.015625,0.015625,0.03125,-0.0078125,0.0,0.015625,0.03125,-0.046875,-0.0234375,0.0390625,-0.015625,0.078125,-0.0859375,-0.0703125,0.046875,0.046875,0.0234375,-0.015625,0.0078125,-0.0859375,-0.0546875,-0.0,0.03125,0.015625,0.0078125,0.0546875,0.0546875,-0.015625,0.0390625,-0.0390625,-0.0078125,0.0078125,0.015625,-0.0078125,0.0,0.015625,-0.0390625,-0.0,-0.0390625,0.015625,0.0078125,-0.0234375,-0.0234375,0.0,-0.015625,0.046875,-0.0234375,0.03125,0.0078125,0.0703125,-0.0078125,-0.0078125,-0.0,0.03125,0.0625,-0.046875,0.078125,0.0078125,0.0078125,-0.015625,-0.0234375,-0.09375,-0.046875,-0.0,0.0,-0.0,0.0078125,-0.0,0.0078125,-0.015625,-0.0,-0.015625,0.0078125,0.03125,-0.078125,-0.0390625,-0.0234375,0.0,-0.0,0.0,-0.0078125,0.0390625,0.03125,-0.03125,-0.0,0.03125,-0.078125,0.015625,-0.0390625,-0.0703125,-0.046875,-0.109375,-0.015625,0.0859375,-0.046875,0.0,-0.015625,-0.0,0.0859375,-0.0234375,0.0390625,0.140625,-0.046875,0.0078125,-0.0703125,-0.0703125,-0.0703125,-0.09375,0.1328125,0.0625,-0.078125,0.0078125,-0.140625,-0.03125,0.1015625,-0.046875,-0.140625,0.046875,-0.0,-0.0234375,-0.015625,-0.0234375,-0.0390625,-0.0859375,-0.0,0.015625,-0.046875,0.0234375,0.0234375,-0.0234375,-0.0234375,0.0,0.015625,0.03125,-0.0078125,0.0625,-0.03125,0.0078125,-0.0,-0.0625,0.046875,0.0078125,0.0390625,0.0546875,-0.0078125,-0.015625,0.015625,0.03125,0.0,-0.0078125,0.046875,-0.03125,0.0859375,-0.0546875,-0.03125,-0.0234375,-0.078125,-0.078125,-0.0234375,0.0078125,0.0703125,0.03125,-0.1015625,-0.0,0.0078125,0.0078125,0.0,-0.015625,-0.015625,-0.0546875,0.046875,-0.015625,0.0703125,0.0703125,-0.03125,-0.0390625,-0.0546875,0.0546875,-0.0234375,0.015625,0.0546875,0.0234375,-0.0078125,0.09375,-0.0625,0.0078125,0.03125,-0.046875,0.109375,0.0390625,0.015625,0.0546875,-0.03125,-0.078125,-0.015625,-0.0546875,-0.0078125,0.0234375,0.0703125,-0.0078125,-0.0546875,0.03125,-0.015625,0.0078125,0.0,0.0859375,0.078125,0.0078125,0.015625,-0.0,0.0078125,0.046875,0.015625,0.0234375,0.0234375,0.03125,-0.0078125,-0.0078125,-0.0,-0.015625,-0.0078125,0.0078125,-0.0,0.015625,0.015625,-0.015625,0.0234375,0.0234375,-0.0078125,0.0546875,-0.0,0.0078125,-0.03125,-0.0234375,-0.0234375,-0.015625,0.0078125,0.0078125,0.015625,0.03125,0.0078125,0.0078125,-0.0,-0.015625,-0.015625,-0.0625,0.015625,-0.046875,-0.0390625,0.0,0.0390625,-0.015625,-0.015625,-0.0,-0.015625,-0.0,0.015625,-0.0078125,-0.0078125,0.0,-0.0078125,0.015625,-0.0390625,-0.015625,0.015625,-0.015625,0.0,0.015625,-0.046875,0.078125,-0.0546875,-0.03125,-0.0078125,0.03125,0.0390625,-0.0078125,-0.0078125,0.0703125,-0.0546875,-0.03125,-0.015625,-0.0234375,0.015625,0.015625,-0.0078125,-0.046875,-0.0390625,0.015625,-0.015625,-0.015625,-0.015625,0.0390625,0.046875,-0.0234375,-0.0,-0.0,-0.0234375,0.03125,-0.015625,0.015625,-0.015625,0.0234375,0.0078125,-0.0078125,0.0546875,-0.015625,0.0,-0.015625,0.015625,-0.0234375,-0.03125,0.03125,0.015625,-0.0234375,0.03125,-0.0,-0.0078125,-0.0078125,0.015625,0.0078125,-0.015625,0.0078125,-0.0,-0.015625,-0.0078125,0.0,0.0234375,-0.015625,-0.0390625,-0.015625,-0.0390625,-0.03125,-0.0078125,-0.015625,-0.0234375,-0.03125,-0.03125,0.0078125,-0.0,-0.03125,0.0625,0.0234375,-0.0078125,-0.03125,-0.0390625,0.0,-0.015625,-0.015625,-0.03125,-0.0,0.0078125,0.0078125,-0.0078125,0.0078125,0.0078125,-0.0078125,-0.015625,0.0078125,0.0078125,-0.015625,-0.0078125,0.015625,0.0390625,0.015625,0.0078125,0.0,0.0703125,0.0078125,0.0078125,-0.0,-0.0234375,-0.03125,0.0390625,-0.078125,-0.03125,-0.0234375,-0.03125,-0.03125,-0.0078125,-0.015625,-0.03125,0.0234375,-0.0625,-0.0546875,0.03125,0.0234375,0.015625,0.03125,-0.03125,-0.046875,-0.015625,-0.1015625,-0.0078125,-0.0234375,0.046875,0.0,0.0,0.015625,0.015625,-0.015625,-0.015625,-0.0546875,0.0546875,-0.0234375,0.0078125,0.0234375,0.015625,0.0078125,0.015625,-0.0234375,0.078125,-0.015625,-0.0234375,0.0234375,-0.015625,0.0234375,-0.0,0.046875,-0.0546875,0.015625,0.0234375,-0.078125,-0.03125,0.0,0.0078125,0.0078125,-0.03125,0.0078125,-0.015625,0.0234375,-0.0234375,-0.015625,0.0078125,0.0078125,0.0625,0.015625,0.0625,0.0859375,-0.03125,-0.015625,-0.03125,-0.046875,-0.0078125,-0.0078125,-0.015625,-0.0546875,-0.03125,0.0234375,-0.0390625,-0.046875,-0.0625,0.0390625,0.0,-0.046875,-0.015625,-0.125,-0.0390625,0.015625,0.0,0.0078125,-0.0390625,-0.03125,0.0078125,-0.1015625,-0.015625,0.0078125,-0.015625,0.0,-0.0234375,0.015625,0.015625,0.0703125,0.0,0.0,-0.015625,-0.03125,-0.03125,0.0546875,-0.0234375,-0.0234375,0.1015625,-0.0078125,0.09375,0.0078125,0.0,-0.015625,-0.0,-0.0078125,0.0078125,0.0390625,0.0078125,-0.0,-0.046875,-0.03125,-0.0078125,0.0390625,0.0546875,0.0078125,-0.0234375,0.0,-0.015625,-0.015625,-0.0390625,-0.015625,0.0078125,-0.0078125,-0.0078125,0.0234375,-0.015625,0.0078125,0.0,-0.0,0.015625,-0.0234375,0.09375,0.109375,-0.0703125,-0.0859375,0.03125,-0.0234375,-0.0078125,-0.0234375,-0.0546875,-0.1328125,-0.0390625,0.0390625,-0.0390625,0.0703125,-0.03125,0.0859375,-0.046875,-0.03125,0.0234375,-0.0546875,0.0625,0.0546875,-0.046875,0.0234375,-0.015625,-0.0625,0.0234375,-0.0078125,0.0078125,-0.0078125,-0.0,-0.0,0.0,-0.0,0.0,0.03125,0.0625,-0.09375,0.0078125,-0.109375,-0.0078125,-0.0546875,0.015625,-0.0625,0.0234375,-0.0234375,0.0390625,-0.1015625,-0.0546875,0.015625,0.03125,-0.0078125,0.046875,-0.0703125,-0.015625,0.109375,-0.09375,-0.015625,0.109375,-0.09375,-0.015625,-0.0234375,0.015625,0.03125,0.1015625,-0.046875,0.0078125,0.0234375,-0.0078125,0.015625,-0.0078125,-0.0390625,-0.0546875,-0.015625,-0.0078125,0.015625,-0.0703125,-0.0390625,0.03125,-0.015625,0.0,-0.046875,0.0,0.046875,-0.03125,-0.0234375,-0.015625,-0.0234375,0.0859375,0.015625,0.03125,-0.015625,-0.0703125,-0.0390625,0.0703125,0.03125,-0.015625,-0.03125,-0.046875,0.0390625,-0.0078125,-0.03125,-0.0390625,0.03125,0.0234375,0.046875,-0.0234375,-0.0390625,-0.015625,0.015625,0.0,-0.015625,-0.0390625,-0.0703125,0.015625,0.0,-0.03125,-0.03125,0.0546875,-0.046875,-0.046875,0.0390625,0.015625,0.03125,0.0,-0.015625,-0.0078125,-0.015625,-0.0078125,0.0078125,0.0078125,0.015625,-0.015625,0.0078125,-0.0546875,0.0625,-0.015625,0.0390625,-0.0078125,0.0234375,-0.03125,0.015625,-0.03125,-0.046875,0.0,0.0,0.0390625,0.015625,0.046875,-0.0390625,-0.0625,0.015625,0.046875,0.0390625,0.0234375,0.0390625,0.0078125,-0.125,0.078125,0.03125,0.0390625,0.09375,0.0234375,-0.078125,0.0546875,-0.015625,-0.03125,0.0234375,0.015625,0.0234375,0.078125,-0.0,-0.0234375,0.015625,0.0390625,-0.0625,0.109375,0.0234375,0.03125,0.09375,0.0078125,-0.078125,0.0078125,-0.0390625,-0.0625,-0.03125,-0.0390625,0.046875,-0.0546875,0.0234375,-0.1328125,0.0078125,0.140625,-0.015625,-0.0859375,-0.0234375,0.140625,0.03125,0.03125,-0.03125,0.0390625,-0.015625,-0.0703125,0.0234375,-0.078125,0.0546875,-0.03125,-0.0390625,0.0234375,-0.0546875,0.03125,0.03125,-0.0234375,-0.0,-0.015625,-0.0390625,0.0078125,0.0390625,-0.09375,-0.0625,0.0390625,0.015625,-0.0078125,-0.0390625,-0.0546875,0.0625,0.015625,-0.140625,0.0546875,0.046875,0.0234375,0.109375,-0.0703125,-0.0234375,0.078125,-0.0078125,0.015625,0.0859375,-0.0234375,-0.015625,-0.046875,-0.125,0.046875,-0.03125,-0.0625,-0.0546875,0.03125,-0.03125,0.0234375,-0.0078125,-0.03125,0.078125,0.0390625,-0.0546875,0.0703125,-0.078125,-0.015625,-0.03125,0.0078125,0.0546875,0.0234375,0.078125,-0.0546875,-0.0078125,0.0234375,-0.0625,0.0,-0.09375,0.0859375,-0.0234375,-0.046875,-0.015625,-0.0625,-0.0625,-0.03125,-0.015625,-0.0390625,-0.0,-0.015625,-0.0078125,-0.0,0.0078125,0.0078125,-0.0,0.015625,0.0078125,-0.0078125,0.0703125,0.125,0.0234375,-0.0078125,-0.0546875,0.0078125,0.0,-0.0703125,0.03125,-0.046875,0.046875,-0.0703125,0.0,-0.078125,0.0,-0.015625,-0.0625,0.0703125,-0.03125,0.03125,0.0234375,0.0859375,-0.03125,0.0703125,0.0,0.0078125,0.0546875,-0.0078125,0.0,-0.015625,-0.0,0.0078125,0.015625,0.0,0.0078125,-0.0078125,-0.015625,-0.046875,-0.015625,0.0078125,0.015625,-0.046875,0.125,0.1015625,-0.0234375,-0.0546875,-0.0078125,-0.0390625,-0.0,0.015625,0.0,-0.0390625,-0.0546875,0.0078125,0.0,0.015625,0.0546875,-0.046875,-0.109375,0.015625,0.046875,-0.0078125,0.0390625,-0.0078125,0.0078125,0.0234375,0.03125,0.0,0.0078125,0.0390625,0.03125,0.015625,0.0,-0.015625,0.0625,-0.0078125,0.0,-0.03125,0.03125,0.0703125,-0.0390625,0.015625,-0.0546875,-0.0234375,0.0078125,-0.0234375,0.0234375,0.03125,0.015625,-0.03125,-0.0078125,-0.015625,-0.046875,0.0,0.0078125,0.0,-0.0078125,-0.0234375,-0.0,-0.0078125,-0.0234375,-0.0078125,-0.0,0.0078125,0.046875,0.0234375,0.0078125,0.015625,0.0078125,0.015625,0.046875,0.046875,0.1171875,-0.0234375,0.0234375,0.0234375,-0.046875,-0.0390625,0.03125,-0.03125,0.015625,0.0859375,-0.0390625,-0.0,0.03125,-0.0390625,-0.015625,0.0,-0.0078125,-0.0078125,-0.0234375,0.0,0.0,-0.0234375,-0.015625,0.0390625,-0.0234375,-0.03125,-0.0078125,0.015625,0.03125,0.0078125,-0.015625,-0.0078125,-0.0390625,0.0234375,-0.0390625,-0.0625,-0.0390625,0.0234375,0.0078125,0.015625,-0.0,0.0234375,0.0703125,0.0546875,0.015625,-0.0234375,-0.0234375,-0.03125,-0.015625,0.03125,-0.0078125,-0.0234375,-0.0546875,-0.0234375,-0.0546875,-0.0625,-0.015625,0.0,0.0078125,-0.015625,-0.0234375,0.015625,-0.0234375,-0.078125,0.0234375,0.03125,-0.0234375,-0.0,0.046875,0.0078125,0.0078125,-0.0234375,-0.0390625,0.015625,-0.0546875,-0.078125,-0.0625,-0.0,0.046875,-0.03125,0.0234375,0.046875,-0.0234375,-0.0546875,-0.09375,-0.015625,0.0625,-0.03125,0.0625,-0.0390625,-0.046875,-0.0390625,-0.0390625,0.0078125,-0.0234375,-0.0078125,0.0546875,0.0234375,-0.046875,-0.015625,-0.03125,-0.046875,-0.078125,-0.03125,-0.0390625,-0.0078125,-0.046875,0.078125,-0.0390625,0.0390625,0.03125,0.0234375,0.078125,0.09375,0.0234375,0.046875,-0.0546875,0.03125,-0.078125,0.03125,0.046875,-0.078125,0.03125,-0.0390625,-0.03125,0.0703125,-0.03125,0.046875,-0.015625,-0.03125,-0.0703125,-0.0234375,0.0,-0.0546875,0.015625,-0.015625,0.0078125,0.0390625,-0.078125,0.015625,-0.0625,0.0546875,-0.046875,0.0234375,0.0390625,-0.0078125,-0.0234375,-0.0234375,-0.03125,-0.0625,-0.078125,-0.0390625,-0.0078125,-0.0234375,-0.046875,-0.03125,-0.0234375,-0.0234375,-0.0234375,-0.0546875,-0.0390625,-0.015625,0.0,0.03125,-0.0078125,0.09375,-0.0234375,-0.015625,-0.0,0.0234375,0.015625,0.0078125,-0.015625,-0.0,0.015625,-0.0078125,0.0234375,0.0078125,0.0,-0.015625,0.078125,0.0546875,0.03125,-0.0078125,0.0234375,0.015625,0.0078125,-0.0,0.0234375,0.03125,-0.015625,-0.0078125,-0.015625,-0.0546875,-0.0234375,0.0078125,-0.0234375,-0.0234375,-0.0390625,-0.046875,0.109375,-0.0234375,-0.03125,-0.015625,0.0078125,0.0,-0.015625,-0.0,-0.0078125,0.0,-0.0,-0.0078125,0.0,-0.0546875,-0.0078125,0.0546875,0.0234375,-0.0546875,-0.0234375,0.0546875,-0.0234375,-0.0390625,-0.0625,-0.0234375,0.0234375,-0.09375,-0.0,0.09375,-0.046875,0.015625,0.0234375,0.0078125,0.0234375,-0.0703125,-0.1171875,0.0390625,0.1015625,-0.0546875,-0.0390625,0.0078125,0.0078125,-0.046875,-0.046875,0.0078125,0.0,-0.015625,-0.046875,0.015625,-0.0390625,0.0234375,0.0546875,-0.0,0.0390625,-0.0078125,-0.0625,0.015625,-0.0078125,-0.015625,-0.015625,0.015625,-0.0,0.0703125,-0.0234375,0.0625,-0.015625,0.0078125,-0.0234375,-0.0234375,0.0078125,-0.03125,-0.0078125,0.03125,0.03125,-0.015625,-0.015625,0.03125,-0.0078125,0.0,0.015625,0.015625,0.015625,0.046875,-0.0390625,-0.0078125,-0.0078125,0.015625,-0.0,-0.046875,0.0234375,0.0546875,-0.09375,0.0078125,-0.0546875,-0.0703125,-0.0546875,-0.0078125,-0.0,0.015625,-0.0703125,0.046875,0.015625,-0.046875,-0.0078125,-0.0,0.0078125,-0.015625,-0.03125,-0.0078125,0.0,-0.0,0.0078125,0.0078125,-0.0078125,0.0078125,0.03125,0.0078125,-0.015625,0.0,-0.03125,-0.0078125,0.0390625,0.09375,-0.03125,-0.0078125,0.015625,-0.0390625,-0.0390625,0.046875,0.015625,-0.015625,0.0,0.015625,-0.109375,-0.015625,-0.03125,0.015625,0.0859375,-0.015625,-0.0078125,0.0234375,0.03125,-0.0859375,0.171875,-0.0625,-0.0390625,-0.0078125,-0.015625,-0.046875,0.0078125,-0.046875,0.03125,0.046875,-0.0390625,-0.015625,-0.046875,-0.09375,-0.0078125,-0.0234375,-0.0234375,-0.0390625,-0.0703125,0.0078125,0.140625,-0.0,-0.0078125,-0.046875,0.0234375,-0.0,-0.03125,-0.0546875,-0.015625,-0.015625,-0.0546875,0.046875,-0.0234375,-0.0390625,-0.03125,-0.0625,0.046875,-0.0546875,0.0546875,-0.0546875,-0.0078125,0.0078125,0.0,-0.015625,-0.015625,-0.0546875,-0.0234375,0.1015625,-0.0859375,-0.0625,-0.0625,-0.0390625,-0.0078125,0.078125,-0.0390625,-0.0078125,-0.0390625,-0.0546875,-0.0078125,-0.0390625,0.0,-0.015625,0.0234375,-0.0,-0.046875,0.078125,-0.0390625,0.0390625,0.0234375,0.0546875,0.0859375,-0.0546875,0.046875,-0.0859375,0.0078125,-0.078125,-0.046875,0.03125,0.0390625,0.046875,0.0625,-0.1328125,-0.015625,0.015625,-0.015625,-0.015625,-0.03125,-0.0390625,0.046875,-0.046875,-0.03125,0.015625,0.0234375,-0.0,-0.0,-0.015625,0.046875,-0.0,0.0390625,-0.046875,-0.0390625,0.046875,0.0078125,-0.0078125,-0.0625,-0.0546875,-0.0234375,-0.0234375,0.0546875,-0.0,0.0,0.0078125,0.015625,0.0078125,0.0,0.015625,-0.0078125,0.0,-0.0,0.0078125,-0.015625,0.0,-0.046875,-0.03125,0.0546875,0.015625,-0.015625,0.015625,-0.0,-0.0078125,-0.0390625,-0.0,-0.0078125,0.0078125,0.015625,-0.0390625,-0.0,-0.015625,-0.0078125,-0.015625,0.0078125,0.0234375,0.046875,0.0078125,-0.046875,0.03125,-0.0078125,-0.03125,0.03125,0.0078125,-0.0078125,0.0,0.0078125,-0.0078125,-0.0,0.0,0.0,-0.0078125,-0.015625,-0.0390625,0.015625,0.015625,0.0078125,0.0078125,-0.015625,-0.0234375,-0.0234375,0.078125,0.03125,0.015625,-0.0390625,-0.0234375,-0.0234375,-0.015625,-0.015625,0.03125,0.0390625,0.046875,-0.015625,-0.0390625,-0.0078125,-0.0390625,-0.015625,0.0,0.0,0.0234375,-0.0,-0.015625,-0.03125,0.0234375,0.015625,-0.0,-0.0234375,-0.0078125,-0.046875,0.078125,-0.015625,0.03125,0.0078125,-0.0390625,-0.0234375,0.0,0.0234375,-0.0078125,0.0546875,-0.0390625,0.015625,-0.0,0.0,0.0078125,-0.0234375,0.0,0.0078125,-0.0078125,-0.015625,0.015625,0.0078125,-0.0078125,0.0,-0.015625,-0.0,0.0234375,-0.015625,0.015625,-0.015625,-0.0234375,0.0234375,-0.0,-0.0078125,-0.0234375,0.0078125,-0.0078125,-0.046875,-0.0546875,-0.0,-0.015625,0.0234375,0.015625,-0.0078125,-0.03125,-0.015625,-0.0546875,-0.0234375,0.0078125,0.0078125,0.015625,0.0234375,-0.0078125,-0.0078125,0.015625,0.0078125,-0.0,-0.0078125,-0.015625,0.015625,-0.0,0.0,-0.0390625,0.0,0.0078125,0.0234375,0.0234375,0.0234375,-0.015625,-0.015625,-0.015625,0.03125,0.0,0.0625,0.0234375,-0.0703125,-0.0078125,-0.0,-0.015625,-0.0078125,0.0703125,0.1171875,-0.0546875,-0.0390625,-0.0,-0.0546875,-0.0234375,-0.0078125,0.015625,-0.0703125,0.03125,0.0390625,-0.015625,-0.0703125,-0.015625,-0.0078125,-0.0234375,0.0078125,0.015625,0.0234375,-0.0234375,0.0,0.0078125,0.0078125,-0.015625,-0.0390625,0.0078125,-0.0390625,-0.0546875,-0.03125,0.0625,-0.0,-0.0625,-0.0078125,0.015625,-0.03125,0.0625,-0.0,0.0703125,0.0390625,-0.1015625,-0.0234375,-0.0234375,0.0234375,-0.0078125,-0.0390625,0.0546875,-0.0,-0.03125,0.0078125,-0.078125,-0.015625,-0.0234375,-0.03125,-0.0078125,0.046875,-0.03125,0.015625,-0.0625,-0.0078125,-0.0234375,-0.0,-0.03125,0.03125,0.0078125,0.0234375,0.0234375,-0.0,-0.03125,-0.03125,0.0078125,0.03125,0.046875,0.03125,0.0078125,-0.0078125,0.0234375,0.03125,0.0,0.0078125,-0.03125,-0.078125,0.0078125,0.078125,0.0390625,-0.0546875,-0.015625,-0.015625,-0.0234375,-0.0390625,-0.0234375,0.015625,0.0546875,0.0078125,0.03125,-0.0078125,-0.0234375,-0.015625,-0.0546875,0.03125,-0.0390625,-0.046875,0.078125,-0.0546875,-0.0234375,0.0078125,-0.0,-0.0078125,-0.046875,0.0078125,-0.015625,0.0078125,0.0234375,0.0078125,-0.015625,-0.015625,0.0234375,-0.0234375,-0.015625,-0.03125,-0.0234375,-0.03125,0.0,-0.015625,-0.0390625,-0.0234375,0.0078125,-0.015625,-0.0078125,-0.0,0.0078125,-0.0078125,-0.0078125,0.0078125,0.0078125,0.0234375,-0.0234375,0.0,-0.0390625,-0.03125,-0.0390625,0.0,0.0078125,0.0078125,-0.0078125,0.0078125,-0.0,-0.03125,0.015625,-0.0234375,0.0,0.0078125,-0.015625,-0.03125,0.0390625,0.015625,0.0234375,0.046875,-0.015625,-0.0234375,-0.0078125,-0.03125,-0.0,0.0,-0.0078125,0.015625,0.0,0.015625,-0.0,0.0078125,0.0078125,0.015625,0.0078125,0.0234375,0.046875,-0.03125,0.0078125,-0.0234375,-0.0078125,-0.015625,0.046875,0.015625,-0.0234375,-0.046875,-0.0,-0.015625,-0.0078125,-0.0234375,0.0,-0.03125,0.046875,0.03125,-0.015625,0.015625,-0.015625,-0.015625,-0.0234375,-0.0390625,-0.0234375,-0.0390625,-0.0234375,0.0,0.0078125,-0.015625,0.0078125,0.0078125,0.0,0.046875,-0.0078125,-0.0,0.0234375,-0.0703125,0.0078125,0.0234375,-0.0078125,0.0234375,0.0546875,-0.0078125,-0.0,0.0078125,-0.015625,0.015625,0.0,-0.015625,-0.0,0.015625,-0.015625,-0.0078125,-0.0,-0.0078125,-0.0078125,0.0078125,0.0078125,0.015625,0.0234375,-0.03125,-0.0234375,-0.03125,-0.0234375,-0.0078125,0.0,0.0,0.0,0.0703125,-0.0234375,-0.0390625,-0.0078125,-0.03125,-0.0,0.0,-0.0234375,0.0234375,-0.078125,0.015625,0.046875,-0.0078125,0.0234375,0.0078125,-0.015625,-0.0078125,0.0234375,-0.0078125,-0.0078125,0.0078125,-0.0078125,-0.0078125,-0.015625,-0.0078125,-0.015625,-0.0078125,-0.0078125,0.0078125,-0.0234375,0.0078125,-0.0078125,-0.0,-0.0,0.0,0.0078125,0.046875,0.015625,0.015625,-0.0234375,0.0078125,-0.03125,-0.0,0.0078125,0.0,0.1796875,0.0234375,0.03125,-0.09375,-0.0390625,0.0078125,-0.015625,-0.0390625,-0.0234375,0.0234375,0.0546875,0.0078125,-0.046875,-0.0078125,-0.0078125,-0.0234375,0.015625,0.03125,-0.03125,-0.015625,-0.0078125,0.03125,-0.0,0.0,-0.0234375,-0.0234375,0.0234375,0.015625,-0.03125,0.03125,0.0078125,0.015625,-0.015625,-0.015625,-0.0234375,-0.0078125,0.0234375,0.0234375,0.0234375,-0.0546875,-0.0078125,-0.046875,-0.0,0.0078125,-0.0,0.03125,0.015625,-0.015625,0.0078125,-0.046875,-0.0078125,0.015625,-0.015625,-0.0078125,0.015625,0.0390625,-0.0078125,0.0390625,0.0546875,-0.015625,0.0,0.0078125,-0.0078125,0.0078125,0.0078125,-0.015625,-0.015625,0.0,0.0078125,-0.0078125,-0.0234375,-0.0078125,0.0859375,0.0234375,-0.0234375,0.0078125,-0.0625,0.0,-0.0078125,0.0078125,0.0,0.03125,0.0234375,-0.0234375,-0.0390625,0.0,-0.0234375,-0.015625,0.0546875,0.0390625,-0.03125,0.03125,-0.0,-0.046875,-0.046875,-0.0078125,0.0078125,0.0078125,0.046875,0.0078125,-0.0546875,-0.0078125,-0.03125,-0.0078125,0.0078125,-0.015625,0.015625,0.0390625,-0.03125,-0.0625,-0.0,-0.0,0.0,0.0078125,0.0234375,-0.0,-0.0,-0.03125,0.046875,0.0703125,-0.0625,0.0234375,0.0546875,0.03125,-0.0078125,0.0078125,-0.0078125,-0.0078125,0.0,-0.0078125,0.015625,-0.0,0.0078125,0.015625,0.0,-0.0390625,0.0703125,0.03125,-0.0546875,0.0078125,0.0,0.015625,-0.046875,0.0546875,0.0,0.0546875,0.0078125,0.0234375,-0.0,-0.0859375,0.0703125,-0.03125,-0.015625,0.0390625,0.015625,-0.03125,0.03125,0.015625,0.078125,-0.0234375,0.03125,-0.0,-0.0078125,0.0078125,-0.0078125,-0.0078125,-0.015625,0.0,0.0,-0.0078125,0.0078125,-0.0,0.046875,-0.0703125,-0.0078125,-0.015625,-0.0,0.0234375,0.015625,-0.078125,0.0546875,-0.0078125,-0.078125,-0.0234375,0.015625,0.015625,-0.046875,-0.015625,0.015625,0.015625,0.03125,-0.0078125,0.015625,0.03125,-0.0234375,0.0078125,-0.0078125,0.0546875,0.0546875,-0.03125,0.03125,0.0078125,-0.0234375,0.0,0.03125,-0.0625,-0.015625,0.0859375,0.0390625,-0.0390625,-0.0234375,0.078125,0.09375,-0.03125,-0.015625,-0.046875,-0.0078125,-0.0703125,-0.0,0.0390625,0.0234375,-0.03125,0.0078125,-0.0078125,-0.015625,-0.0390625,0.0078125,-0.015625,0.0,-0.0234375,0.0078125,0.0,0.015625,0.0,-0.015625,-0.0390625,0.03125,0.1015625,-0.0546875,0.0,-0.0234375,0.0,0.0078125,0.0,-0.0546875,-0.0,-0.0546875,0.0703125,0.03125,0.03125,-0.0625,-0.0625,-0.015625,0.1015625,-0.03125,-0.03125,0.0078125,0.046875,-0.0390625,-0.0078125,0.0546875,0.0078125,-0.0078125,-0.0078125,0.015625,0.0078125,0.0234375,-0.0,0.0078125,0.0078125,-0.0234375,0.0078125,0.0234375,0.0390625,-0.0390625,0.015625,0.0625,0.015625,0.0,-0.0234375,-0.0703125,0.0078125,0.0078125,-0.03125,-0.0078125,0.0234375,0.03125,-0.046875,0.0078125,-0.09375,-0.0078125,-0.0703125,-0.109375,-0.0,0.0546875,-0.0234375,0.078125,-0.0078125,-0.109375,-0.046875,0.0,-0.015625,0.0078125,-0.0234375,0.0546875,0.0390625,0.0078125,-0.0,0.03125,-0.0390625,-0.0234375,0.0390625,0.0546875,0.015625,-0.015625,-0.0,-0.015625,0.0390625,-0.0078125,-0.0078125,0.0234375,-0.0078125,-0.046875,0.0234375,-0.015625,-0.0234375,0.015625,-0.0546875,-0.109375,-0.0859375,-0.0234375,0.0,0.046875,0.0859375,0.03125,-0.0390625,0.03125,0.0234375,0.015625,0.0078125,-0.0234375,-0.0390625,0.0078125,0.0,-0.0234375,-0.0703125,0.03125,-0.015625,-0.0234375,0.046875,-0.0078125,-0.078125,-0.078125,0.0234375,0.015625,-0.0078125,0.015625,0.0078125,-0.0,0.0078125,0.03125,0.1484375,0.0234375,-0.015625,-0.03125,-0.0546875,-0.03125,-0.03125,-0.0,0.0546875,-0.0546875,-0.015625,0.015625,-0.0703125,-0.0625,-0.0234375,0.0703125,-0.0703125,-0.0859375,0.0703125,0.046875,-0.0703125,-0.0859375,0.03125,0.0546875,-0.0703125,0.0625,0.0078125,-0.0390625,0.0546875,-0.0234375,-0.03125,-0.0625,-0.0078125,0.0390625,-0.0234375,0.0078125,0.0859375,0.0390625,-0.09375,-0.078125,-0.015625,0.015625,-0.078125,0.015625,0.0078125,0.0234375,0.015625,-0.015625,-0.0390625,0.0078125,0.03125,0.0546875,0.0625,0.0,-0.015625,-0.015625,-0.0,-0.0078125,-0.015625,-0.0078125,-0.0078125,-0.0,0.0546875,0.015625,0.0703125,0.0390625,-0.0625,0.0078125,-0.03125,-0.015625,0.0,0.0234375,0.0546875,0.0078125,0.03125,-0.0234375,-0.0,-0.0234375,-0.015625,-0.015625,-0.0,-0.046875,0.0078125,-0.046875,0.03125,-0.015625,0.015625,0.0078125,-0.015625,0.0078125,-0.0078125,-0.0078125,-0.0078125,-0.015625,0.0078125,-0.0078125,0.0078125,0.0078125,0.03125,-0.015625,-0.0,-0.015625,-0.046875,0.015625,0.0078125,-0.03125,-0.0,-0.0234375,-0.046875,-0.0859375,0.0625,0.0390625,-0.015625,0.03125,-0.0078125,0.046875,0.0234375,-0.015625,-0.0234375,-0.0703125,-0.0078125,-0.015625,-0.0546875,-0.0625,-0.015625,0.015625,0.015625,-0.015625,0.078125,-0.0,0.0078125,-0.0,0.0,0.015625,0.0234375,0.0390625,-0.0234375,-0.03125,0.015625,-0.03125,-0.0078125,-0.046875,-0.0234375,-0.0078125,-0.0234375,-0.0234375,0.0078125,-0.0078125,-0.0078125,0.015625,-0.0078125,0.0078125,0.0,0.0078125,-0.0078125,-0.015625,-0.0078125,-0.015625,-0.0234375,0.0078125,0.046875,0.0234375,-0.0,0.03125,0.0390625,-0.046875,0.0078125,-0.015625,-0.015625,-0.0234375,0.0,-0.03125,-0.0078125,0.0625,0.0390625,-0.0078125,0.03125,-0.0390625,-0.015625,-0.015625,-0.03125,0.0234375,0.0078125,-0.0234375,-0.015625,0.0390625,0.0234375,-0.046875,-0.0078125,-0.0,-0.0078125,-0.0,-0.015625,0.015625,-0.015625,-0.015625,-0.0078125,0.0,-0.0234375,-0.015625,0.0078125,0.0,-0.015625,0.0,0.0078125,0.03125,0.0078125,0.03125,0.0078125,0.046875,0.03125,-0.03125,0.0234375,0.015625,0.0234375,0.0234375,-0.03125,-0.03125,0.03125,0.03125,-0.03125,0.0,-0.0546875,-0.0234375,-0.015625,0.0078125,-0.0078125,-0.0,0.03125,0.0546875,-0.0234375,-0.03125,-0.015625,0.015625,-0.03125,-0.03125,0.0234375,0.03125,-0.015625,-0.0078125,-0.0078125,0.0234375,0.0078125,-0.0078125,0.0078125,0.0078125,-0.015625,0.0078125,-0.0078125,0.0078125,0.015625,0.015625,0.0078125,0.1015625,-0.03125,-0.0625,-0.0234375,-0.03125,0.0234375,0.03125,-0.03125,-0.0234375,0.0078125,-0.0,-0.0390625,-0.015625,0.0078125,0.015625,0.0078125,0.0078125,-0.015625,0.0078125,0.0,0.015625,-0.0,-0.0234375,-0.0546875,0.0078125,-0.0,-0.015625,-0.0234375,-0.03125,-0.0078125,-0.0078125,-0.015625,0.0078125,-0.0078125,-0.0234375,-0.0390625,0.015625,0.046875,-0.0546875,0.046875,-0.0078125,-0.046875,-0.03125,-0.03125,-0.0234375,-0.03125,-0.015625,0.0703125,-0.015625,0.015625,-0.0234375,-0.015625,0.0390625,0.0390625,0.0703125,0.015625,-0.0,-0.015625,-0.0390625,-0.0546875,0.0078125,-0.0078125,-0.0703125,0.015625,0.0,-0.0078125,0.0234375,0.015625,0.0078125,0.03125,0.0078125,0.03125,-0.0078125,-0.03125,-0.0234375,-0.0703125,0.0078125,0.0390625,0.0625,-0.09375,0.0546875,0.015625,-0.0078125,0.0390625,0.015625,0.078125,0.09375,-0.0,0.0078125,-0.0078125,0.0078125,0.0234375,-0.0,-0.015625,0.015625,-0.0078125,-0.0078125,0.0234375,-0.0234375,0.03125,0.0546875,-0.0390625,-0.03125,0.0078125,-0.015625,0.0,0.0078125,-0.015625,-0.015625,0.0078125,-0.0234375,-0.0234375,-0.03125,-0.0546875,0.0078125,0.0234375,-0.0078125,-0.0078125,0.0234375,-0.015625,0.0234375,-0.0390625,-0.0546875,0.0,0.0,-0.0,0.015625,-0.015625,-0.015625,-0.0,0.0,-0.0078125,0.0078125,-0.0546875,0.015625,-0.015625,0.015625,-0.0,-0.0234375,-0.046875,-0.0625,0.0,0.0234375,0.0234375,-0.0234375,-0.0234375,-0.0078125,0.0703125,0.0078125,-0.0546875,0.046875,0.0625,-0.0,0.0078125,-0.0859375,-0.0078125,-0.0078125,-0.0546875,-0.0390625,-0.0078125,0.0078125,-0.0625,0.0078125,0.0078125,0.0625,-0.0390625,0.0078125,0.0390625,0.015625,-0.0703125,0.0703125,0.015625,-0.0,-0.0625,0.0078125,-0.0390625,-0.03125,0.0234375,-0.0078125,0.03125,-0.03125,-0.0,-0.0078125,0.0,-0.015625,-0.03125,0.0,-0.015625,-0.015625,-0.0078125,0.015625,-0.0234375,0.0078125,0.015625,0.0,0.0078125,0.046875,-0.0390625,0.0078125,-0.015625,-0.0546875,-0.0234375,-0.015625,-0.046875,0.0078125,0.0078125,0.015625,0.015625,-0.078125,-0.0390625,0.0078125,0.0390625,0.1015625,0.0859375,-0.0859375,0.0234375,-0.0234375,-0.0234375,-0.03125,-0.0078125,-0.015625,0.0,0.0234375,-0.0078125,0.0078125,-0.0,-0.015625,0.0,0.0,-0.0,0.015625,-0.0078125,-0.0078125,0.015625,-0.015625,-0.0,0.0625,-0.046875,-0.015625,-0.03125,-0.03125,0.03125,-0.0078125,-0.0078125,-0.0234375,-0.0703125,-0.046875,-0.0,0.0,-0.0390625,0.140625,0.015625,-0.0,-0.1171875,-0.078125,-0.046875,-0.0703125,-0.03125,-0.0,-0.078125,-0.0234375,0.0390625,-0.078125,-0.09375,-0.0,0.046875,-0.0390625,0.0078125,-0.0,0.0078125,-0.03125,0.0625,0.0546875,-0.046875,0.015625,-0.0078125,-0.0,-0.0390625,0.0,-0.0390625,-0.015625,0.0390625,-0.03125,0.0234375,-0.0,0.0,0.15625,-0.0625,-0.046875,-0.0,-0.1015625,-0.0234375,-0.0546875,-0.0546875,-0.0625,-0.03125,-0.0,-0.0234375,-0.0390625,-0.0234375,-0.046875,-0.0,-0.015625,-0.0078125,-0.0703125,-0.0546875,-0.015625,-0.015625,-0.015625,-0.046875,-0.0078125,-0.0078125,-0.0234375,0.078125,-0.0078125,-0.0078125,0.015625,0.0,-0.0078125,-0.0546875,-0.0390625,0.0234375,0.0078125,-0.0078125,-0.0234375,-0.03125,-0.0078125,0.0,-0.0390625,-0.0234375,0.0625,-0.0078125,-0.046875,0.015625,-0.03125,-0.046875,0.046875,-0.03125,-0.03125,0.078125,0.015625,-0.015625,-0.015625,0.03125,0.03125,-0.0390625,-0.03125,-0.1015625,0.0234375,0.0,-0.0,-0.015625,0.0703125,-0.0078125,0.0,0.0546875,-0.0078125,0.0234375,-0.078125,0.0078125,-0.0,0.078125,0.0078125,0.0078125,-0.015625,-0.046875,0.0234375,-0.0234375,-0.046875,-0.0703125,0.0078125,-0.0078125,-0.0390625,0.0,0.0546875,-0.0234375,0.0078125,0.0078125,-0.0078125,0.015625,-0.015625,0.015625,0.015625,0.0078125,0.0078125,-0.0,-0.03125,-0.0,-0.0625,-0.0234375,0.0390625,0.03125,0.015625,0.0,0.015625,-0.0234375,-0.0,0.0,-0.0234375,-0.0078125,0.0078125,-0.0390625,-0.0546875,-0.0390625,0.09375,-0.0078125,0.015625,-0.0078125,-0.0234375,0.0390625,-0.0078125,0.0078125,0.0078125,0.0078125,-0.0,0.0,0.0078125,-0.0,0.0078125,0.015625,0.0,0.03125,-0.0390625,-0.015625,-0.0078125,-0.03125,0.0546875,0.03125,0.0,0.0703125,-0.046875,-0.046875,0.0859375,-0.0390625,-0.0390625,0.0390625,0.015625,-0.1015625,0.0234375,-0.046875,0.0625,-0.0078125,-0.0390625,-0.0546875,-0.109375,-0.0078125,0.0390625,-0.03125,-0.0,0.03125,-0.0078125,-0.0078125,0.015625,-0.0,0.0,0.015625,-0.046875,-0.015625,0.0546875,-0.0390625,-0.0390625,-0.046875,-0.046875,-0.0078125,0.0859375,0.0546875,0.0234375,0.0234375,0.03125,0.0234375,-0.015625,0.015625,0.03125,0.015625,-0.015625,0.0390625,0.015625,0.046875,-0.0234375,-0.03125,0.015625,-0.0,-0.015625,-0.0078125,-0.0,-0.0078125,0.03125,0.0078125,-0.0546875,-0.046875,0.0078125,-0.0390625,-0.0625,-0.0,-0.0,-0.140625,-0.0390625,-0.0546875,0.0234375,-0.03125,0.046875,-0.0234375,-0.0390625,-0.0078125,0.109375,0.015625,-0.046875,-0.0703125,0.015625,0.0546875,0.0390625,0.0078125,0.015625,0.0078125,-0.0078125,0.0078125,-0.0,-0.0078125,0.0,-0.0078125,0.0625,0.015625,0.03125,0.0,0.015625,-0.015625,0.0234375,-0.0234375,-0.0234375,0.0078125,0.015625,-0.03125,-0.0078125,-0.0859375,0.046875,0.0078125,0.0234375,0.015625,-0.03125,-0.03125,-0.0078125,-0.0234375,-0.0703125,0.2421875,0.0234375,0.0390625,-0.1171875,-0.0234375,-0.0,0.0078125,-0.0234375,-0.0625,-0.015625,-0.0234375,-0.0390625,0.0078125,-0.0,0.0546875,-0.0,-0.03125,-0.0078125,-0.1015625,0.015625,0.0703125,0.0234375,-0.0,-0.0,0.0078125,-0.0078125,-0.03125,-0.046875,0.0390625,0.078125,0.0078125,0.0390625,-0.03125,0.0234375,-0.0078125,-0.046875,0.046875,0.0078125,0.015625,-0.0546875,-0.0234375,0.03125,-0.0,-0.0,0.0625,-0.0234375,0.015625,-0.0078125,-0.0390625,-0.015625,-0.046875,-0.0078125,-0.015625,0.015625,-0.046875,-0.015625,0.078125,0.09375,0.03125,-0.015625,0.0234375,-0.0234375,-0.0234375,-0.0390625,0.0703125,0.0234375,0.0390625,-0.015625,0.03125,0.015625,-0.0625,-0.0234375,-0.03125,-0.0078125,-0.0,0.046875,-0.0,0.046875,-0.0390625,-0.0234375,0.015625,0.0703125,-0.0390625,-0.0546875,-0.0859375,-0.0234375,-0.0390625,-0.078125,-0.0625,-0.03125,0.0,-0.046875,0.015625,0.0234375,-0.0390625,0.078125,0.0859375,-0.0234375,-0.03125,0.09375,-0.0078125,0.03125,0.015625,0.03125,-0.0625,-0.0078125,-0.0234375,-0.0390625,-0.03125,-0.0234375,0.078125,0.0859375,0.0078125,0.0546875,-0.0390625,0.015625,0.015625,0.0,-0.0546875,-0.0078125,-0.0234375,-0.0078125,-0.0,0.0,-0.0,-0.0,-0.0078125,-0.0078125,0.0078125,0.0078125,0.0234375,0.0703125,0.0546875,-0.03125,-0.046875,-0.015625,0.046875,0.0859375,0.0234375,-0.0234375,-0.0390625,-0.0078125,-0.015625,-0.0546875,0.109375,0.015625,0.046875,-0.0234375,0.0078125,-0.0,0.0390625,0.0390625,-0.015625,0.0234375,-0.0078125,-0.078125,-0.03125,-0.0078125,-0.0078125,-0.0,0.015625,-0.0078125,0.0078125,0.0078125,-0.0078125,-0.0078125,-0.0,-0.046875,-0.078125,-0.0703125,0.0078125,-0.015625,0.0546875,0.0859375,-0.03125,0.0234375,-0.0390625,-0.046875,-0.015625,0.0078125,0.0078125,0.0234375,-0.046875,-0.015625,-0.0390625,-0.03125,-0.0390625,-0.015625,0.0078125,0.0546875,-0.046875,0.0078125,-0.03125,0.0,-0.0,0.0390625,-0.03125,-0.09375,-0.0234375,0.0390625,0.046875,-0.015625,-0.0234375,-0.03125,-0.015625,0.015625,0.0390625,0.0078125,-0.0078125,0.0390625,-0.0078125,-0.03125,-0.0546875,0.0546875,0.0,-0.015625,0.0078125,-0.015625,-0.03125,0.0390625,0.03125,-0.015625,-0.0078125,0.0,0.03125,-0.03125,0.0,-0.0234375,0.0078125,0.015625,0.03125,-0.015625,-0.03125,-0.0078125,0.015625,0.0,-0.0625,-0.046875,0.0234375,-0.0234375,-0.0546875,0.0390625,0.03125,0.078125,-0.046875,-0.0078125,-0.0625,-0.0390625,0.0546875,0.015625,0.03125,-0.0078125,-0.046875,0.0234375,-0.0078125,-0.0390625,0.0078125,0.0078125,0.0,0.0,-0.0,-0.0,0.0234375,0.0,-0.0,0.015625,-0.03125,-0.0,-0.0078125,-0.03125,-0.015625,0.0546875,0.0234375,-0.0078125,0.0625,-0.1328125,0.03125,0.0390625,0.03125,0.0078125,0.015625,-0.03125,-0.03125,0.03125,-0.0078125,-0.0546875,0.046875,-0.0546875,0.0625,-0.0,0.015625,0.0,0.078125,0.0234375,0.0078125,-0.03125,-0.0390625,-0.0703125,0.0078125,0.015625,-0.0390625,0.0234375,-0.0078125,0.0546875,-0.0234375,-0.0546875,0.03125,0.0625,-0.0546875,0.0234375,0.0234375,-0.03125,-0.0078125,0.0,-0.03125,-0.0078125,-0.03125,0.03125,0.0078125,0.0625,-0.0625,0.03125,0.0703125,-0.0625,-0.015625,0.09375,-0.0078125,0.0390625,-0.03125,0.0234375,0.0234375,-0.0390625,0.0078125,0.0,0.0390625,0.015625,0.046875,-0.03125,-0.0078125,0.109375,0.03125,0.0078125,0.046875,0.03125,-0.0078125,0.0234375,-0.03125,0.0234375,0.0390625,-0.0546875,0.046875,-0.015625,-0.0234375,-0.046875,0.015625,0.046875,0.0546875,-0.0234375,-0.0625,0.0078125,-0.046875,0.046875,-0.0546875,-0.0,0.0078125,-0.0,-0.0234375,-0.0078125,0.078125,0.0078125,0.0078125,-0.0546875,-0.0078125,0.0390625,-0.0546875,0.0078125,-0.046875,-0.0390625,-0.0546875,0.03125,0.0078125,0.0390625,-0.015625,0.03125,-0.046875,-0.0234375,0.0390625,-0.0390625,-0.03125,0.0078125,0.0078125,0.1171875,-0.09375,-0.015625,0.0625,-0.046875,-0.0234375,0.0234375,0.0,0.015625,0.03125,-0.09375,-0.0546875,-0.046875,0.0078125,-0.0078125,0.03125,-0.015625,-0.0390625,0.0078125,0.0078125,0.0,-0.015625,-0.0,0.0,0.0,0.015625,0.0,0.0234375,-0.0,-0.0,-0.0,0.0078125,-0.078125,-0.0625,0.0078125,-0.0234375,-0.03125,0.015625,0.0,-0.0,-0.0625,-0.015625,0.0078125,-0.0,0.0078125,0.0625,0.0390625,0.0234375,0.046875,0.03125,-0.015625,-0.0234375,-0.046875,-0.0078125,0.015625,-0.015625,0.0078125,0.0,0.0,0.0078125,0.0078125,-0.0078125,-0.0,-0.015625,-0.0078125,0.015625,-0.0078125,-0.125,0.078125,0.0078125,0.0703125,-0.09375,0.015625,0.0546875,-0.015625,0.0703125,0.046875,0.0,-0.046875,0.03125,0.0546875,0.015625,0.0390625,0.0390625,-0.0234375,-0.0,-0.09375,0.0234375,-0.0,0.015625,-0.0234375,0.0,-0.0,-0.015625,0.046875,-0.09375,-0.0,-0.015625,0.015625,-0.03125,0.03125,-0.0078125,0.046875,-0.0234375,0.046875,0.0625,-0.0078125,-0.03125,0.03125,-0.015625,-0.0234375,-0.0546875,0.0390625,-0.0078125,-0.03125,-0.015625,0.0234375,-0.0078125,0.0390625,-0.015625,-0.015625,-0.015625,-0.0078125,-0.03125,0.015625,0.0390625,0.0625,0.0234375,-0.0234375,-0.0390625,-0.0390625,-0.03125,0.0234375,0.03125,-0.0078125,-0.078125,-0.0625,0.0,-0.0234375,-0.0390625,0.0078125,0.0703125,0.0234375,-0.015625,-0.015625,-0.0078125,0.0,0.109375,-0.046875,-0.046875,-0.046875,-0.015625,-0.0703125,0.0,-0.0078125,-0.0,0.015625,-0.0,-0.015625,-0.0,-0.015625,-0.0078125,-0.0,-0.015625,-0.015625,-0.0390625,0.0078125,-0.015625,-0.0,-0.015625,-0.0625,-0.0078125,-0.0234375,-0.0078125,-0.0234375,0.078125,-0.0078125,0.015625,-0.0390625,0.0078125,-0.0234375,0.046875,0.0078125,-0.0078125,-0.0,-0.0234375,-0.0078125,-0.015625,-0.0234375,0.0234375,-0.0703125,-0.015625,-0.0078125,0.03125,0.0078125,0.015625,0.0,-0.015625,0.0390625,-0.03125,-0.0390625,-0.0546875,-0.0,-0.0390625,0.0703125,-0.0625,0.015625,0.09375,-0.0078125,0.015625,-0.015625,-0.0390625,-0.0390625,-0.0078125,-0.046875,0.015625,-0.0390625,0.046875,0.015625,-0.0078125,-0.0546875,0.0859375,-0.0703125,0.0078125,0.0078125,-0.0078125,0.0,-0.0234375,-0.046875,0.0390625,-0.0625,0.0234375,0.0546875,-0.015625,-0.015625,-0.0078125,0.0078125,-0.03125,0.0234375,-0.0078125,-0.0546875,0.125,0.1015625,0.046875,0.078125,-0.046875,-0.0078125,-0.0546875,-0.0546875,-0.03125,0.015625,0.0625,-0.0390625,0.0078125,-0.0078125,0.1015625,-0.125,-0.0390625,0.0234375,0.0078125,-0.015625,-0.0078125,-0.0234375,0.03125,0.0859375,0.0546875,0.0546875,-0.03125,-0.0234375,-0.046875,0.015625,0.0390625,0.03125,-0.015625,-0.0234375,-0.03125,-0.015625,0.1171875,0.015625,0.03125,0.0703125,0.0625,0.0234375,-0.03125,-0.0234375,-0.046875,-0.0234375,-0.0390625,0.0078125,0.0078125,0.0234375,-0.0078125,-0.015625,0.0625,0.0,-0.0234375,-0.0078125,-0.0078125,0.0234375,0.0078125,0.0234375,-0.0546875,0.140625,-0.0,-0.046875,0.0078125,-0.0078125,0.015625,-0.0078125,-0.0,0.03125,0.0,-0.0078125,0.0234375,-0.0,-0.015625,-0.0,0.078125,-0.1015625,0.015625,0.0390625,-0.0703125,-0.0078125,-0.03125,-0.0546875,-0.0546875,0.015625,0.0,-0.0390625,0.0234375,-0.0234375,0.015625,0.0,-0.0546875,-0.0,-0.0390625,-0.046875,0.03125,0.0078125,0.0,-0.0625,0.03125,0.015625,-0.015625,-0.0078125,-0.015625,-0.0078125,-0.0,0.0078125,-0.0,0.0078125,0.1171875,0.0703125,0.0859375,-0.03125,-0.15625,0.0546875,0.0234375,-0.0390625,-0.0,-0.03125,-0.0390625,-0.03125,0.1015625,0.015625,-0.0390625,-0.0234375,-0.0703125,0.046875,-0.03125,0.1328125,-0.0390625,-0.0390625,0.0859375,-0.140625,-0.046875,-0.046875,-0.078125,0.03125,-0.03125,0.0078125,-0.0078125,-0.03125,-0.0,0.0234375,-0.0546875,-0.0234375,0.046875,0.125,-0.0078125,-0.046875,-0.015625,0.0,-0.015625,0.0,-0.0,0.0078125,-0.03125,0.03125,0.046875,-0.03125,0.0,0.03125,-0.0078125,0.03125,0.0,-0.0546875,-0.0,-0.0,-0.0,-0.046875,0.0,-0.0078125,0.0234375,-0.015625,-0.0078125,-0.0546875,-0.03125,0.0234375,-0.0234375,0.0234375,0.03125,-0.0078125,-0.015625,0.0546875,0.015625,-0.0703125,0.046875,0.0234375,-0.078125,-0.1015625,0.0078125,-0.0703125,0.0234375,0.0703125,-0.0625,0.0625,-0.0078125,-0.0234375,0.015625,-0.046875,-0.0078125,0.0078125,0.0078125,-0.015625,-0.0078125,0.015625,-0.0078125,0.0,-0.015625,-0.0234375,-0.046875,0.0234375,-0.0,-0.0390625,0.0,-0.0,-0.046875,0.046875,0.0390625,-0.1171875,-0.046875,0.015625,-0.015625,-0.0078125,-0.0703125,-0.015625,0.015625,-0.015625,0.0859375,-0.0546875,-0.0078125,0.0390625,0.015625,0.015625,-0.03125,0.0234375,-0.0625,0.1015625,0.0078125,-0.0390625,-0.0546875,-0.0,-0.0078125,-0.046875,0.0859375,-0.0625,-0.0625,-0.0078125,-0.0546875,-0.0625,-0.0078125,-0.0390625,-0.0078125,-0.046875,0.015625,-0.03125,0.078125,0.078125,-0.0078125,-0.0078125,-0.0234375,-0.015625,-0.078125,-0.140625,0.046875,-0.015625,-0.046875,0.0859375,-0.078125,-0.015625,-0.03125,-0.0078125,-0.0703125,0.0390625,-0.046875,-0.0546875,0.015625,-0.125,-0.015625,0.09375,0.015625,-0.0625,0.0390625,-0.0546875,-0.03125,-0.0078125,-0.03125,-0.0625,0.0390625,-0.0234375,0.0078125,-0.0625,-0.0625,0.0234375,0.015625,0.0234375,-0.0390625,-0.0390625,-0.03125,0.0078125,0.03125,0.046875,-0.0390625,0.0,-0.0,-0.03125,0.0546875,-0.0546875,-0.0390625,0.015625,0.09375,-0.046875,-0.0546875,-0.1171875,0.03125,0.1015625,0.109375,-0.0234375,0.0625,0.046875,-0.0546875,-0.0390625,-0.0078125,-0.03125,0.015625,-0.046875,-0.0234375,-0.0625,0.0625,-0.03125,0.0078125,-0.0,0.0234375,0.0234375,0.109375,0.15625,-0.0546875,0.0234375,0.0390625,-0.03125,0.0390625,-0.0234375,0.0078125,-0.0,0.046875,-0.0390625,-0.0390625,-0.03125,0.0546875,-0.046875,0.109375,0.0078125,0.0625,0.0078125,-0.0078125,0.015625,-0.0078125,0.0078125,-0.015625,0.0,0.0078125,0.015625,0.0078125,0.0625,0.0078125,-0.0859375,-0.0,-0.03125,0.0546875,-0.046875,-0.0078125,-0.0390625,-0.0703125,0.0078125,-0.0234375,-0.015625,-0.0234375,0.0703125,-0.0625,-0.0703125,-0.0078125,-0.0078125,-0.046875,0.0625,-0.0234375,-0.046875,-0.0234375,0.03125,-0.015625,0.0078125,-0.0078125,-0.015625,-0.0078125,0.0,0.0078125,-0.0078125,-0.0078125,-0.0078125,0.0,0.0546875,0.015625,-0.0234375,-0.046875,-0.078125,-0.0546875,-0.125,-0.0234375,0.015625,0.09375,-0.078125,0.0,-0.015625,-0.0390625,-0.0,0.015625,0.0,-0.1015625,-0.0625,-0.0625,0.0078125,0.0,-0.0,0.0625,-0.0078125,-0.0390625,0.0234375,-0.03125,0.0390625,0.0234375,-0.0234375,-0.0859375,0.015625,0.046875,-0.0234375,-0.0390625,0.046875,-0.0078125,-0.0703125,0.015625,0.0234375,0.0234375,-0.0546875,0.0234375,-0.078125,-0.046875,-0.03125,0.0078125,0.0,0.0078125,-0.0234375,0.0078125,0.015625,-0.0546875,0.0,0.0078125,-0.0234375,-0.0234375,0.03125,0.015625,-0.015625,0.0,-0.0234375,-0.0234375,0.0,-0.0546875,-0.015625,-0.015625,-0.0625,-0.03125,-0.046875,0.0078125,0.0,-0.03125,0.046875,0.015625,0.0546875,0.171875,-0.0703125,0.015625,0.015625,0.0625,0.0,-0.0390625,-0.0234375,-0.0234375,0.1328125,0.03125,-0.015625,-0.0078125,-0.0078125,0.0078125,0.015625,-0.015625,0.0078125,0.0,-0.03125,0.0,-0.0,-0.015625,0.0,-0.0234375,0.03125,-0.046875,-0.0,-0.0703125,0.0078125,-0.0703125,-0.046875,-0.0703125,-0.03125,0.0625,-0.0078125,-0.0625,0.0078125,-0.046875,-0.046875,0.0390625,-0.03125,-0.0546875,-0.03125,-0.0078125,0.0390625,-0.0625,0.0703125,0.0078125,-0.015625,-0.015625,0.046875,-0.0234375,-0.0703125,-0.03125,-0.0234375,-0.046875,-0.03125,-0.0390625,0.0234375,-0.078125,0.03125,0.0078125,0.0625,0.171875,0.0078125,-0.0390625,0.0703125,-0.03125,-0.03125,0.1484375,-0.0390625,-0.0546875,-0.03125,0.015625,0.03125,-0.078125,-0.046875,-0.1015625,0.1015625,0.03125,-0.0703125,-0.015625,-0.0625,0.0234375,-0.0234375,0.03125,-0.015625,-0.015625,0.0078125,-0.0234375,-0.0390625,0.0078125,-0.0625,-0.046875,-0.046875,0.015625,-0.0625,0.0,-0.0625,-0.015625,-0.0625,-0.078125,-0.0390625,-0.0234375,0.015625,0.046875,0.03125,-0.015625,-0.0078125,-0.078125,0.0234375,-0.0390625,-0.03125,0.0078125,-0.09375,0.0625,-0.0546875,-0.046875,-0.015625,-0.046875,0.03125,-0.0625,0.0,0.03125,0.0234375,0.09375,0.03125,-0.046875,-0.046875,0.03125,-0.0234375,-0.046875,-0.1015625,0.0,-0.046875,0.0,0.0078125,-0.0546875,0.1796875,-0.03125,-0.0859375,0.09375,0.0,0.0,-0.109375,-0.0546875,-0.0234375,-0.0703125,-0.0078125,-0.0703125,0.0625,-0.015625,-0.015625,0.0,-0.03125,0.0234375,-0.046875,-0.0078125,-0.0546875,0.0546875,0.015625,-0.0234375,-0.0390625,0.0390625,0.0078125,0.0,0.0078125,0.015625,-0.015625,-0.0078125,0.0,-0.0,-0.0078125,0.03125,-0.046875,-0.0390625,0.015625,-0.0078125,0.03125,-0.0078125,-0.015625,-0.015625,0.0,0.0078125,-0.03125,0.0,-0.0078125,0.0234375,0.0,-0.0078125,-0.0546875,0.03125,0.03125,-0.0390625,-0.0546875,0.015625,0.078125,-0.0234375,0.0,0.015625,-0.0,-0.0078125,-0.0078125,0.0078125,0.0078125,0.0078125,0.0078125,-0.0078125,0.015625,0.03125,-0.0,-0.0,0.046875,-0.0078125,-0.015625,0.015625,-0.0546875,-0.0234375,-0.0078125,-0.0390625,0.0,-0.0234375,0.0390625,-0.03125,-0.0625,-0.03125,-0.03125,-0.0390625,-0.015625,0.0078125,-0.0859375,-0.0,0.0703125,-0.015625,0.015625,-0.0546875,0.03125,-0.03125,0.015625,-0.0390625,-0.0390625,-0.0078125,-0.0,-0.0078125,-0.0078125,-0.015625,-0.0625,-0.0546875,0.0390625,-0.0390625,-0.015625,0.0234375,0.0078125,0.03125,-0.0,-0.0078125,-0.015625,-0.0078125,-0.0234375,0.015625,-0.015625,-0.0078125,-0.0078125,0.0078125,-0.0078125,-0.0078125,-0.0078125,-0.0078125,-0.015625,-0.015625,-0.03125,-0.0,-0.046875,-0.0078125,-0.03125,-0.03125,-0.0390625,0.046875,-0.0078125,0.0078125,-0.015625,0.0390625,0.0078125,-0.046875,0.0390625,0.0,-0.015625,0.015625,0.0234375,0.0234375,0.015625,-0.0078125,0.078125,-0.0234375,0.015625,0.0234375,0.0234375,0.0078125,0.0,0.015625,0.015625,0.0,-0.0078125,0.015625,0.03125,-0.0,-0.0078125,-0.0078125,-0.03125,-0.0,-0.0390625,0.0,0.0234375,-0.0390625,0.0234375,0.015625,0.0390625,0.0078125,0.0234375,0.015625,0.046875,-0.0234375,-0.0234375,-0.046875,-0.0546875,-0.03125,0.046875,-0.0078125,-0.015625,0.0234375,0.015625,0.03125,0.015625,-0.0234375,-0.0546875,0.046875,-0.0,-0.0078125,0.015625,0.03125,-0.0625,-0.03125,-0.03125,-0.0234375,0.0078125,-0.0078125,-0.0078125,-0.0546875,-0.0390625,0.0234375,-0.015625,-0.015625,-0.0,0.078125,0.015625,-0.0234375,0.0546875,-0.015625,0.0,0.015625,0.015625,-0.03125,-0.03125,-0.0,0.046875,0.078125,0.0078125,-0.0625,-0.0234375,-0.0078125,-0.0546875,-0.03125,0.0234375,-0.09375,-0.0234375,0.046875,0.0390625,-0.0078125,0.0859375,0.0625,-0.0,0.0,-0.0234375,-0.0390625,-0.0,0.03125,-0.015625,0.015625,0.046875,0.03125,0.0390625,-0.015625,0.015625,0.1015625,0.0390625,-0.03125,-0.0390625,-0.0234375,-0.1015625,-0.046875,0.1015625,-0.0234375,-0.0078125,0.0390625,0.0234375,-0.03125,-0.0546875,0.0078125,-0.078125,-0.046875,0.046875,0.078125,-0.0625,-0.03125,-0.046875,0.015625,-0.03125,-0.1015625,-0.0390625,0.0078125,-0.0703125,0.0234375,-0.015625,-0.046875,-0.0,0.015625,0.03125,-0.046875,0.03125,-0.0234375,-0.0390625,0.0078125,0.0,-0.0078125,-0.078125,-0.046875,-0.0,-0.03125,-0.03125,0.0390625,0.0078125,-0.0078125,-0.015625,0.015625,-0.0,-0.046875,0.0625,0.0546875,-0.03125,-0.0390625,-0.0078125,0.0,-0.0078125,0.015625,0.015625,-0.0,0.015625,-0.0,-0.015625,-0.015625,0.0,0.0390625,-0.0234375,-0.0,0.0546875,-0.0234375,0.0078125,-0.0234375,0.015625,0.015625,0.046875,0.015625,0.0078125,0.015625,-0.015625,-0.0546875,-0.0234375,-0.015625,0.078125,-0.03125,0.03125,0.0390625,-0.0078125,0.046875,-0.0078125,-0.015625,-0.0234375,-0.0,0.0078125,-0.0078125,0.0078125,-0.0,-0.0078125,-0.0078125,-0.0078125,-0.0078125,0.0078125,-0.015625,-0.0,-0.03125,0.0,-0.046875,0.015625,-0.03125,-0.0,0.0546875,0.0,-0.03125,-0.0625,0.109375,-0.015625,-0.0078125,-0.0625,0.0078125,0.0234375,0.03125,-0.015625,0.015625,-0.0078125,-0.0390625,0.015625,-0.0625,-0.0078125,0.03125,0.0,-0.0234375,-0.0078125,0.0,-0.046875,0.0625,0.0234375,0.03125,0.0078125,0.0078125,0.0078125,-0.03125,-0.03125,0.0078125,0.046875,-0.0390625,-0.015625,0.015625,-0.0078125,-0.015625,-0.015625,-0.046875,-0.046875,0.015625,-0.0,-0.0234375,-0.03125,0.0078125,-0.0,-0.0234375,0.03125,0.0078125,-0.0390625,-0.0,-0.015625,0.0,-0.0,0.015625,-0.015625,0.015625,-0.0078125,0.0078125,-0.0234375,-0.03125,-0.0078125,-0.0546875,-0.03125,0.0234375,-0.03125,-0.0078125,0.0703125,-0.015625,-0.03125,0.015625,-0.046875,-0.0390625,0.0703125,-0.03125,-0.03125,0.046875,-0.0234375,-0.03125,-0.0625,0.0078125,-0.015625,0.0078125,-0.0,-0.0078125,0.0,0.0078125,-0.0,-0.0,-0.015625,0.0078125,0.03125,-0.03125,-0.015625,-0.03125,-0.0,0.0234375,0.03125,-0.046875,-0.0234375,0.0625,0.0625,-0.015625,-0.0546875,0.03125,-0.015625,-0.0078125,-0.015625,-0.046875,-0.015625,0.0234375,0.0546875,0.0390625,-0.0078125,-0.0078125,0.09375,-0.0234375,-0.0,0.078125,0.015625,-0.0234375,-0.0703125,-0.0,-0.0390625,-0.0546875,-0.0234375,0.015625,0.0234375,0.015625,0.046875,0.0390625,-0.0625,-0.046875,-0.015625,0.0390625,0.0,-0.046875,0.046875,0.0234375,-0.03125,-0.046875,-0.0234375,-0.0234375,-0.03125,-0.0390625,0.0546875,0.03125,-0.0546875,-0.0859375,0.03125,0.0234375,-0.0625,0.03125,0.0234375,-0.03125,-0.0078125,0.0078125,-0.0,-0.0078125,0.015625,0.015625,0.0234375,0.015625,-0.0078125,-0.0078125,-0.0078125,0.046875,-0.03125,-0.0546875,-0.0390625,0.0078125,0.0078125,0.03125,-0.03125,0.03125,0.0078125,-0.0234375,-0.0390625,0.0078125,-0.03125,-0.0703125,0.0390625,-0.046875,-0.03125,0.0703125,-0.015625,-0.046875,-0.03125,0.0,-0.015625,0.03125,0.015625,-0.0,-0.046875,0.0625,0.0,0.03125,0.0234375,-0.015625,0.0390625,0.0546875,-0.046875,-0.0234375,-0.0234375,-0.015625,-0.0078125,0.0078125,0.0234375,-0.015625,0.0546875,0.0078125,-0.0625,0.0,0.015625,0.0078125,0.015625,0.046875,0.0546875,0.03125,-0.0234375,-0.0390625,-0.0234375,0.0,-0.0,-0.0390625,0.015625,-0.0234375,-0.0078125,0.0078125,-0.0546875,0.0078125,0.0,-0.03125,-0.0,-0.015625,-0.0,-0.0078125,-0.0,0.0234375,0.015625,-0.0078125,-0.0,0.0859375,0.015625,-0.0078125,0.0234375,0.0,-0.0078125,0.03125,0.0234375,-0.0078125,0.078125,0.015625,-0.03125,0.046875,0.015625,-0.0078125,-0.0078125,0.0390625,0.0078125,-0.03125,-0.03125,-0.015625,-0.015625,0.046875,-0.0078125,-0.0,-0.0546875,-0.0234375,-0.0078125,-0.0078125,0.0,0.0078125,0.0078125,0.0078125,0.0078125,0.0078125,-0.0078125,0.015625,0.1015625,0.015625,-0.046875,-0.0546875,-0.0078125,-0.0546875,0.0078125,-0.0390625,0.0546875,-0.0546875,0.03125,-0.0390625,0.046875,-0.0,-0.0078125,-0.03125,-0.0546875,-0.03125,-0.0234375,0.0234375,-0.0625,0.1328125,0.0078125,-0.015625,0.046875,-0.0078125,0.0,0.015625,-0.0078125,0.03125,-0.015625,-0.0,0.0,-0.0390625,-0.015625,0.0234375,-0.0078125,0.03125,-0.0859375,0.0390625,0.078125,-0.015625,-0.0234375,-0.0078125,0.0,-0.0390625,-0.03125,0.0390625,-0.015625,-0.0390625,-0.0,-0.0078125,0.046875,0.03125,0.0390625,0.03125,0.0,-0.0,0.03125,-0.0234375,-0.0078125,0.0390625,0.0234375,-0.0078125,-0.03125,0.015625,-0.0625,-0.0234375,-0.0078125,0.0078125,-0.0,-0.03125,-0.0625,0.015625,-0.0078125,-0.0078125,-0.0546875,0.0078125,0.0078125,0.046875,-0.0625,-0.0625,0.0234375,-0.0,0.0859375,0.03125,-0.0,-0.0390625,-0.046875,0.0078125,-0.0,-0.0,-0.0078125,-0.015625,0.0078125,-0.0078125,0.0,0.0,0.078125,-0.015625,-0.03125,-0.0234375,-0.0234375,-0.0234375,0.0078125,-0.0078125,-0.015625,-0.0234375,0.0,-0.0390625,-0.015625,-0.0,-0.015625,0.0390625,0.0703125,-0.03125,-0.0703125,-0.046875,0.125,0.0078125,-0.046875,-0.1015625,0.0546875,-0.0546875,-0.0078125,0.046875,-0.0,-0.0390625,-0.0390625,-0.0546875,0.0546875,-0.03125,0.015625,-0.03125,0.015625,0.0625,0.0078125,0.0625,-0.0703125,-0.015625,0.015625,-0.0703125,-0.0078125,0.0,0.0234375,-0.0234375,-0.015625,0.0390625,-0.0390625,0.015625,0.0390625,-0.0,0.03125,-0.0390625,0.046875,0.015625,0.0,-0.046875,-0.03125,0.046875,-0.0078125,-0.0078125,-0.046875,-0.0078125,-0.03125,-0.0234375,-0.0234375,0.0390625,0.0546875,0.0703125,-0.015625,-0.0078125,-0.0390625,-0.03125,-0.015625,0.03125,0.015625,0.03125,-0.0078125,0.046875,-0.0234375,0.0390625,0.03125,-0.0546875,-0.0234375,0.015625,-0.0546875,0.0078125,0.0390625,-0.078125,-0.0390625,-0.0,-0.03125,-0.0703125,-0.0078125,0.0234375,-0.0,0.015625,0.03125,-0.0390625,-0.0390625,-0.015625,0.0078125,-0.03125,0.0234375,0.0078125,0.09375,0.03125,-0.0,-0.0,-0.0625,0.03125,-0.03125,-0.0078125,0.0078125,0.0390625,0.0,0.03125,-0.0078125,-0.046875,0.0625,0.0234375,0.0,-0.0234375,-0.0234375,-0.0234375,0.0,-0.0546875,0.0,-0.0390625,-0.046875,0.0234375,0.015625,-0.0,-0.0625,-0.0078125,-0.0078125,0.015625,0.0234375,0.0234375,-0.0390625,-0.015625,-0.015625,-0.0078125,-0.0,-0.0078125,0.0,0.015625,-0.0,0.0078125,-0.0078125,0.0078125,0.0625,0.0078125,0.0546875,-0.015625,-0.015625,0.015625,-0.0390625,0.0078125,0.0234375,-0.0703125,0.03125,0.0234375,0.1015625,-0.046875,0.0078125,-0.015625,-0.0546875,0.078125,0.0703125,-0.0234375,-0.0703125,-0.0703125,0.0078125,-0.0546875,-0.0078125,-0.0078125,0.015625,0.0,-0.0,0.0078125,-0.0078125,0.0,-0.0078125,0.0078125,0.0,-0.0078125,-0.015625,0.046875,0.0390625,-0.0234375,-0.0546875,0.0078125,-0.0,-0.015625,-0.0625,-0.015625,-0.0625,0.0390625,0.046875,0.0390625,0.09375,-0.03125,0.015625,-0.0234375,-0.0546875,0.015625,0.03125,0.0234375,0.015625,-0.03125,-0.0625,-0.0234375,-0.0078125,-0.0078125,0.0078125,-0.0078125,-0.0390625,-0.0078125,0.0390625,-0.0,0.0078125,0.0078125,0.0078125,0.0078125,-0.03125,0.0,0.015625,-0.0703125,-0.0390625,0.0078125,-0.015625,-0.0078125,-0.03125,-0.0078125,-0.015625,-0.0078125,-0.015625,-0.015625,-0.0078125,-0.0234375,-0.0,-0.0390625,0.0078125,-0.015625,-0.015625,0.0,-0.0078125,0.015625,0.0234375,-0.0390625,-0.03125,0.0078125,-0.03125,0.0,-0.0078125,-0.0078125,-0.03125,-0.0078125,-0.0546875,0.0390625,-0.0,0.0,0.0078125,0.0859375,-0.0078125,-0.0234375,0.0546875,0.015625,-0.0078125,-0.046875,0.0078125,0.0546875,-0.0390625,-0.015625,-0.0234375,0.015625,0.015625,0.0078125,-0.0,-0.0078125,-0.0,-0.0078125,-0.015625,-0.0078125,0.03125,0.0,0.03125,-0.0078125,0.0078125,-0.015625,0.0234375,-0.03125,0.0546875,-0.03125,-0.0078125,-0.046875,-0.03125,0.046875,-0.0625,-0.015625,0.015625,-0.0234375,-0.046875,-0.0078125,0.0234375,0.03125,-0.0625,-0.0703125,0.0078125,-0.015625,0.0234375,0.0,-0.0390625,-0.0234375,-0.0078125,-0.0,-0.0078125,-0.015625,-0.0234375,-0.03125,-0.0,0.1015625,-0.03125,-0.046875,-0.0859375,-0.015625,-0.0078125,0.0234375,0.0390625,0.0078125,-0.015625,0.0078125,-0.0078125,0.0625,-0.046875,-0.0234375,0.046875,-0.0390625,-0.0234375,0.0546875,-0.0078125,-0.046875,-0.03125,-0.0390625,-0.0078125,-0.0,-0.078125,0.0859375,0.0,-0.0234375,-0.0390625,-0.015625,-0.0625,-0.0546875,0.0,0.03125,-0.0234375,0.0,-0.015625,-0.03125,0.046875,0.015625,-0.046875,0.078125,0.0546875,-0.015625,-0.0078125,-0.0390625,0.015625,0.0859375,-0.0234375,-0.015625,-0.0625,0.0234375,-0.03125,0.0078125,0.0703125,-0.0078125,-0.09375,0.0390625,-0.0078125,-0.0625,0.0,0.0625,-0.0234375,0.046875,0.0546875,-0.0234375,-0.0078125,-0.0625,0.015625,-0.0078125,-0.046875,0.03125,-0.0078125,0.0078125,0.0390625,-0.015625,-0.015625,-0.0390625,-0.015625,-0.046875,-0.015625,0.03125,-0.0078125,0.03125,-0.03125,0.03125,0.0078125,-0.0234375,-0.0234375,0.0234375,-0.0078125,-0.0390625,-0.0078125,-0.03125,-0.0078125,0.078125,-0.015625,-0.0703125,-0.0234375,-0.0078125,-0.046875,0.015625,0.015625,-0.0234375,-0.0078125,0.0234375,0.015625,0.0,0.0078125,0.015625,-0.0078125,-0.015625,-0.0078125,0.0078125,0.015625,0.0546875,-0.015625,0.015625,0.015625,0.015625,0.03125,-0.015625,-0.015625,-0.03125,0.0078125,0.046875,0.046875,-0.0390625,-0.0078125,-0.015625,-0.015625,0.015625,-0.015625,0.0078125,0.0078125,-0.046875,0.046875,-0.015625,-0.0078125,0.0,-0.015625,-0.0234375,0.0078125,0.0,-0.0078125,0.0078125,-0.0,0.0078125,-0.0,-0.0078125,-0.015625,-0.03125,0.015625,-0.015625,0.046875,0.046875,-0.03125,-0.015625,-0.0234375,-0.015625,0.125,-0.03125,-0.015625,-0.078125,-0.03125,-0.03125,-0.0078125,-0.0234375,0.0078125,-0.0234375,0.0078125,0.03125,-0.0625,-0.0078125,-0.0546875,-0.0078125,-0.03125,-0.015625,0.015625,-0.0078125,0.0,0.0078125,0.015625,0.0,-0.0078125,-0.0234375,0.015625,-0.0078125,0.0078125,-0.0078125,0.0234375,-0.0234375,-0.03125,-0.03125,-0.015625,0.015625,0.0078125,0.0234375,-0.0078125,0.0390625,-0.0390625,-0.0078125,0.0078125,-0.0234375,-0.0078125,0.0078125,-0.015625,-0.015625,-0.0078125,-0.0,0.0,0.0078125,-0.0078125,0.015625,0.0078125,0.015625,-0.0,-0.078125,-0.015625,0.0,0.015625,0.0,0.0,0.125,-0.046875,-0.03125,-0.1015625,-0.046875,-0.03125,-0.0078125,-0.0,-0.0,-0.0859375,0.0546875,-0.0546875,-0.03125,-0.0078125,-0.0,-0.0078125,0.0078125,0.0390625,-0.0234375,-0.015625,0.015625,-0.0,-0.0078125,-0.0078125,0.0078125,0.0,-0.0078125,-0.0234375,0.0078125,-0.0078125,-0.015625,0.03125,0.03125,-0.015625,-0.0,-0.0078125,0.0625,-0.078125,0.015625,0.0078125,0.015625,0.0078125,-0.03125,0.0234375,0.03125,0.2890625,0.0703125,-0.0390625,-0.1875,-0.046875,-0.0625,-0.0390625,-0.0078125,-0.0078125,0.03125,-0.0390625,-0.015625,-0.03125,0.015625,0.0234375,-0.03125,-0.0078125,0.0078125,-0.0390625,-0.0234375,-0.015625,0.03125,-0.0078125,0.0390625,-0.0390625,-0.0625,0.0,-0.015625,-0.0625,0.0,0.0078125,0.046875,0.0703125,-0.0078125,-0.0,0.0078125,0.1015625,-0.015625,0.0390625,-0.03125,-0.0859375,0.0,-0.015625,-0.0078125,-0.0,0.0390625,0.0234375,-0.0078125,0.015625,-0.0859375,-0.0234375,-0.0234375,-0.0390625,0.015625,-0.0078125,-0.0390625,0.0234375,0.03125,0.03125,0.046875,0.015625,0.0,-0.0234375,-0.0078125,0.0078125,-0.03125,-0.0546875,-0.015625,-0.0546875,0.015625,-0.0078125,-0.015625,0.0703125,-0.0078125,-0.03125,-0.046875,-0.0390625,-0.0,-0.015625,0.03125,-0.03125,0.1015625,-0.0390625,0.0078125,-0.0234375,-0.0625,-0.0078125,-0.0234375,-0.015625,0.03125,0.03125,0.03125,0.0234375,0.015625,0.015625,0.0234375,-0.0234375,-0.046875,-0.015625,0.015625,-0.0625,-0.0234375,0.03125,-0.0234375,0.0546875,-0.0234375,0.015625,0.015625,-0.0234375,-0.046875,-0.015625,-0.015625,-0.046875,0.03125,-0.0234375,-0.0078125,0.0234375,-0.015625,-0.0390625,0.0078125,0.125,-0.0078125,-0.0234375,-0.0234375,0.03125,-0.0078125,-0.015625,-0.0078125,0.0078125,0.015625,0.0,-0.0,0.015625,-0.0,0.0078125,-0.0,0.0234375,-0.0078125,0.03125,-0.0859375,-0.046875,-0.0234375,-0.0078125,-0.0234375,-0.03125,-0.015625,0.0390625,-0.0234375,0.0625,0.03125,0.0,0.0078125,-0.015625,-0.0390625,0.046875,-0.0078125,-0.0390625,0.0,0.015625,0.1171875,0.0390625,-0.015625,0.0,0.0078125,-0.0078125,0.0,-0.0078125,-0.0,-0.0078125,-0.0078125,0.0078125,-0.015625,-0.0,-0.03125,-0.0234375,-0.0703125,-0.015625,0.0,-0.0625,-0.0390625,0.0234375,0.0234375,-0.0078125,0.0078125,0.0625,-0.0078125,0.0234375,0.0234375,-0.015625,-0.09375,-0.046875,0.078125,0.03125,-0.0390625,0.015625,0.0546875,-0.015625,-0.0234375,0.0625,-0.0078125,-0.0234375,0.046875,0.0078125,-0.0546875,-0.0546875,0.015625,-0.0234375,0.015625,-0.0234375,-0.0390625,0.0625,0.0,-0.015625,0.0390625,-0.0078125,-0.015625,0.03125,-0.03125,-0.0234375,0.046875,0.0234375,0.0390625,-0.03125,-0.015625,0.0078125,-0.03125,0.0234375,-0.0078125,-0.015625,-0.0078125,0.015625,0.0078125,0.0234375,0.015625,0.0078125,0.0078125,-0.0,0.0234375,-0.015625,0.03125,0.015625,-0.0703125,-0.0234375,-0.0234375,-0.0703125,-0.0390625,0.0,0.0546875,-0.046875,0.0078125,0.0078125,-0.015625,-0.03125,-0.03125,-0.03125,-0.125,-0.0078125,0.0078125,0.0703125,0.09375,-0.0078125,-0.0078125,-0.0078125,-0.0078125,-0.015625,-0.0,0.0078125,0.03125,0.03125,-0.0078125,0.03125,0.0390625,0.0,0.0078125,-0.046875,-0.0,0.0078125,0.0234375,-0.0078125,0.0,-0.0078125,-0.0234375,-0.0390625,0.0546875,-0.015625,0.015625,0.0546875,-0.015625,-0.03125,-0.0390625,-0.0234375,-0.1015625,-0.046875,-0.0390625,0.0546875,0.0078125,-0.0078125,0.0078125,-0.078125,-0.0390625,-0.0390625,-0.0390625,0.0078125,0.1015625,0.0859375,-0.0234375,0.03125,0.0703125,-0.0390625,-0.109375,0.0,-0.015625,-0.0234375,0.0390625,-0.046875,-0.0703125,0.03125,0.0234375,0.046875,-0.0078125,-0.03125,0.015625,-0.015625,-0.0,0.015625,-0.0078125,-0.015625,-0.015625,-0.015625,-0.0234375,0.0390625,-0.1015625,-0.0234375,0.03125,-0.03125,-0.0,-0.046875,-0.03125,-0.015625,-0.0234375,-0.0078125,-0.0234375,0.0390625,-0.015625,0.0,0.0703125,-0.0078125,0.0390625,-0.0703125,-0.0390625,-0.0234375,0.0234375,0.0078125,-0.0234375,-0.0390625,0.0859375,-0.0078125,0.078125,0.0625,-0.0078125,-0.140625,0.0703125,0.0,-0.1328125,-0.046875,0.0234375,0.03125,-0.1328125,-0.03125,0.046875,-0.015625,-0.046875,-0.0078125,-0.03125,-0.0234375,-0.015625,-0.0546875,-0.0234375,0.1015625,0.0234375,-0.0078125,0.0078125,0.0234375,0.0078125,-0.015625,-0.0546875,-0.015625,-0.0078125,0.015625,-0.0078125,0.0859375,-0.0546875,0.0078125,-0.0078125,-0.0390625,0.0,0.046875,0.0390625,-0.0234375,-0.03125,-0.015625,0.0078125,-0.03125,-0.0546875,-0.0,-0.0546875,0.0859375,-0.0546875,-0.0234375,-0.0546875,-0.03125,0.0234375,0.0859375,0.0234375,0.015625,0.0,-0.0234375,0.0,-0.0078125,-0.015625,0.015625,0.015625,-0.0,-0.0859375,0.046875,-0.0703125,0.046875,-0.03125,-0.03125,0.0234375,0.078125,-0.0234375,-0.0,-0.0234375,-0.0,0.0390625,-0.015625,-0.0078125,0.0078125,-0.0234375,0.0234375,-0.03125,-0.078125,-0.015625,0.0078125,-0.015625,0.0078125,0.0234375,0.03125,-0.0234375,-0.0078125,0.015625,-0.0078125,-0.0,-0.0078125,-0.015625,0.0,0.0078125,0.0078125,-0.0625,-0.0234375,-0.03125,-0.015625,-0.046875,0.0078125,0.0078125,-0.015625,0.0234375,-0.0546875,0.0390625,0.0,0.0,-0.0390625,-0.03125,-0.0390625,-0.015625,-0.03125,-0.0078125,-0.015625,-0.015625,0.03125,0.015625,0.0390625,-0.015625,-0.046875,-0.0078125,-0.0625,-0.0078125,0.0078125,0.0,0.0078125,0.03125,-0.0390625,-0.015625,-0.0078125,0.0,-0.0078125,-0.015625,-0.0703125,0.0234375,-0.03125,-0.0234375,-0.0390625,-0.0234375,-0.03125,-0.0078125,-0.0234375,0.0234375,-0.0234375,-0.0078125,-0.0,0.0078125,-0.0234375,0.0078125,0.0078125,0.0390625,-0.0078125,0.0,-0.0,-0.015625,-0.0078125,-0.0,-0.0078125,-0.0234375,0.0,0.078125,0.0078125,-0.0078125,-0.0234375,-0.0078125,-0.0390625,-0.015625,-0.046875,-0.0234375,-0.03125,0.0078125,-0.0390625,-0.015625,-0.015625,0.015625,0.03125,0.0546875,-0.0625,0.0078125,-0.0390625,-0.015625,0.015625,0.0390625,-0.0,-0.0078125,-0.015625,0.0078125,0.015625,0.0234375,0.046875,-0.0,0.0,0.0078125,-0.0234375,0.0390625,0.0078125,0.015625,-0.0234375,0.0078125,0.0234375,-0.0234375,-0.046875,0.0546875,-0.0390625,0.078125,-0.0,-0.0,-0.0234375,-0.015625,-0.0078125,0.0078125,-0.03125,-0.046875,-0.03125,-0.0390625,-0.03125,-0.03125,-0.03125,0.0078125,0.0078125,-0.0,-0.078125,0.046875,0.0234375,-0.0234375,-0.015625,0.0390625,0.0390625,0.0078125,0.0234375,-0.0,-0.0078125,0.0078125,-0.0546875,0.0078125,-0.0,-0.03125,-0.03125,-0.09375,-0.0078125,-0.03125,-0.0078125,-0.0,-0.0390625,0.0234375,0.03125,0.0546875,0.0234375,0.0078125,0.078125,-0.015625,-0.015625,-0.0078125,-0.03125,-0.0078125,-0.0234375,-0.0078125,0.0625,-0.0390625,-0.0078125,-0.0234375,-0.0390625,0.03125,0.015625,0.0078125,-0.0,0.0859375,0.03125,0.0,-0.0234375,0.015625,0.03125,-0.0703125,0.0234375,0.015625,-0.03125,0.0078125,0.0,0.046875,0.078125,-0.0390625,0.0546875,-0.0546875,0.0546875,0.03125,0.0390625,0.015625,-0.0078125,-0.0390625,0.0078125,0.0234375,-0.03125,0.09375,-0.0703125,-0.015625,-0.0,0.09375,0.078125,0.0234375,-0.0390625,0.015625,-0.015625,0.0234375,0.0078125,0.0078125,0.0,0.0859375,0.0390625,-0.046875,-0.0390625,-0.0625,0.046875,-0.0234375,-0.03125,-0.0703125,-0.0546875,0.0703125,0.0390625,0.03125,0.0234375,0.0546875,0.0234375,-0.0546875,-0.109375,-0.0390625,-0.0234375,-0.015625,-0.0234375,0.0625,0.0390625,-0.0859375,-0.0390625,-0.0234375,0.046875,-0.03125,0.015625,0.0703125,0.0,-0.0078125,0.03125,0.015625,-0.0234375,-0.0234375,0.015625,0.0078125,0.0078125,0.03125,0.0078125,-0.03125,-0.015625,-0.03125,-0.0078125,-0.0078125,-0.0234375,0.0390625,-0.0078125,0.078125,-0.0,-0.0390625,0.0078125,-0.0078125,-0.0234375,-0.0546875,-0.0078125,0.0078125,-0.0390625,-0.109375,0.0546875,0.0234375,-0.0234375,-0.0234375,-0.0625,0.03125,-0.015625,-0.0078125,-0.0,-0.0,-0.0,-0.0,-0.0078125,0.0078125,-0.0,0.0234375,0.0625,0.0234375,-0.046875,-0.03125,-0.0625,0.03125,-0.0546875,-0.015625,0.03125,-0.0546875,-0.015625,0.0703125,-0.0078125,-0.0546875,-0.046875,-0.0859375,0.0234375,0.1015625,-0.0625,-0.03125,-0.078125,-0.09375,0.0390625,-0.015625,-0.015625,0.1171875,0.0,0.0078125,0.0,0.0,0.0078125,-0.0625,0.0078125,-0.03125,0.015625,0.0390625,0.0703125,0.046875,-0.0078125,0.125,-0.015625,-0.0546875,-0.0078125,-0.015625,-0.0,-0.015625,0.0234375,-0.0390625,-0.0625,0.015625,0.03125,-0.0234375,-0.0078125,-0.03125,-0.0234375,0.0078125,0.0234375,0.0390625,-0.03125,0.0,-0.015625,-0.03125,-0.015625,0.0,0.0390625,0.046875,-0.0703125,-0.0,0.0078125,0.0078125,0.0,-0.0546875,-0.03125,-0.03125,0.0078125,0.0703125,0.0078125,-0.0703125,-0.03125,0.0078125,0.0859375,0.0234375,-0.015625,-0.078125,0.046875,-0.0078125,-0.03125,-0.0078125,0.0234375,0.0234375,0.0234375,-0.0,0.0,-0.0,0.0,-0.0078125,0.0,-0.0,0.0390625,0.015625,-0.046875,-0.03125,0.0390625,-0.015625,0.0,-0.0234375,-0.0234375,-0.1015625,-0.078125,0.0390625,0.0,-0.09375,0.015625,0.0078125,-0.0,-0.0078125,-0.015625,0.046875,0.0078125,-0.0390625,-0.046875,0.0078125,-0.0078125,-0.0546875,0.0546875,0.078125,0.0234375,0.015625,-0.0390625,-0.0390625,-0.0703125,-0.03125,-0.0234375,-0.0546875,-0.0390625,0.0546875,-0.046875,-0.046875,0.015625,-0.0078125,-0.03125,-0.078125,-0.0390625,-0.0078125,0.109375,-0.0390625,0.0,-0.1328125,0.0078125,-0.015625,0.0390625,-0.0078125,-0.03125,-0.078125,-0.0390625,0.1171875,-0.0859375,0.0234375,0.03125,-0.015625,0.015625,-0.0078125,-0.015625,0.0078125,0.0,0.046875,0.0078125,-0.046875,-0.0390625,-0.0078125,-0.046875,0.0390625,0.015625,0.0078125,-0.046875,-0.0078125,-0.046875,-0.09375,0.0234375,-0.0234375,-0.046875,-0.0234375,0.0546875,0.0078125,-0.046875,0.0234375,-0.0390625,0.0078125,-0.078125,-0.03125,0.0234375,-0.0703125,0.046875,0.0703125,-0.0625,0.1015625,-0.0078125,-0.0625,-0.03125,0.0234375,0.046875,-0.015625,-0.046875,0.015625,-0.0078125,-0.015625,-0.0546875,-0.0,0.0625,0.1015625,0.15625,-0.046875,-0.0078125,-0.03125,-0.0234375,0.109375,0.015625,0.0625,0.109375,-0.0078125,-0.015625,0.015625,0.015625,-0.0078125,-0.0078125,0.1015625,-0.0546875,-0.03125,0.015625,0.0625,-0.0,-0.0703125,-0.0234375,-0.0390625,-0.0859375,0.0078125,-0.0625,-0.0234375,-0.0,-0.046875,-0.03125,-0.046875,-0.0078125,-0.0,-0.0078125,-0.0078125,-0.015625,0.0078125,0.0078125,0.0078125,0.0078125,0.046875,0.0859375,0.0390625,-0.0078125,0.09375,-0.1328125,-0.0625,0.015625,-0.0625,0.0,-0.0234375,0.015625,-0.0234375,0.0234375,-0.015625,-0.015625,-0.0234375,-0.109375,-0.0234375,0.0390625,-0.0078125,0.0078125,-0.0703125,0.1171875,0.0078125,-0.0625,-0.046875,-0.0078125,-0.0,-0.015625,0.015625,-0.015625,0.015625,-0.015625,-0.015625,0.0078125,-0.015625,-0.0234375,-0.0625,-0.046875,0.0546875,0.03125,-0.0234375,-0.046875,-0.0625,0.09375,-0.0703125,0.03125,-0.0390625,-0.1171875,-0.0546875,-0.046875,0.0078125,-0.03125,0.0078125,0.140625,-0.0078125,-0.15625,0.0703125,-0.1640625,0.046875,-0.0234375,-0.015625,-0.0078125,0.0390625,-0.0234375,0.0,0.0546875,-0.0703125,-0.0234375,0.0,-0.0546875,-0.0,0.0625,-0.03125,0.0234375,-0.0234375,-0.0078125,-0.0234375,0.0,0.046875,0.0,-0.0234375,0.0078125,-0.0234375,0.0078125,0.03125,0.0078125,0.046875,-0.015625,0.0859375,0.0390625,0.015625,-0.0,0.0390625,-0.015625,-0.0234375,-0.0234375,0.03125,-0.0,0.0625,0.015625,0.015625,0.0078125,0.015625,-0.03125,0.015625,-0.0390625,-0.046875,-0.0703125,0.078125,-0.03125,-0.0390625,-0.03125,-0.0078125,-0.1015625,0.046875,-0.046875,0.0390625,-0.0625,-0.0390625,-0.0078125,0.046875,-0.03125,-0.0703125,0.0546875,-0.0078125,-0.0078125,-0.0078125,-0.0078125,-0.015625,-0.0234375,0.0078125,-0.015625,-0.0078125,-0.0078125,-0.1328125,0.0078125,-0.0078125,0.0078125,-0.0078125,-0.0234375,0.0078125,-0.0390625,0.0703125,-0.0703125,0.0703125,-0.015625,-0.0078125,-0.046875,0.0,0.078125,-0.046875,0.0234375,-0.0390625,-0.0,-0.03125,-0.0546875,-0.03125,0.03125,-0.0625,0.0390625,0.046875,-0.03125,0.03125,0.03125,0.015625,-0.03125,-0.03125,-0.0859375,-0.0625,-0.0078125,-0.09375,0.0390625,-0.078125,-0.046875,0.046875,-0.0859375,0.0078125,0.1640625,0.015625,-0.0078125,-0.0625,-0.046875,0.09375,-0.0078125,-0.0390625,-0.0234375,-0.0625,-0.0390625,-0.1015625,-0.0234375,0.1640625,0.09375,0.015625,-0.1171875,0.1484375,-0.0859375,0.015625,-0.03125,0.046875,0.0390625,0.0546875,0.015625,-0.0859375,-0.0078125,0.0078125,-0.0078125,-0.015625,-0.03125,-0.03125,-0.0078125,-0.0078125,-0.125,-0.0234375,-0.03125,0.0390625,0.09375,0.0625,0.015625,-0.0625,-0.03125,0.03125,0.03125,0.125,-0.015625,0.0234375,0.0078125,0.0546875,0.0390625,-0.03125,-0.0703125,0.03125,0.0234375,-0.0390625,-0.0625,-0.015625,0.0390625,0.0,0.0234375,-0.0546875,0.015625,0.03125,0.0078125,0.015625,0.0234375,0.015625,0.03125,0.0234375,-0.0625,0.0546875,-0.03125,0.0,-0.03125,-0.015625,-0.0546875,0.015625,-0.0234375,-0.03125,-0.015625,-0.0390625,0.0234375,-0.1328125,0.0,-0.015625,-0.0703125,-0.046875,-0.015625,0.15625,-0.0,0.0234375,0.0390625,0.0078125,0.0078125,-0.0390625,-0.0234375,0.078125,0.03125,-0.0234375,0.0234375,-0.0,-0.0078125,0.0078125,-0.0078125,0.0078125,-0.0078125,-0.0,0.0234375,-0.015625,0.0234375,0.0234375,-0.03125,-0.0390625,-0.0390625,0.0546875,-0.046875,-0.0234375,-0.0078125,-0.0546875,-0.0078125,-0.046875,0.0234375,-0.0078125,0.0234375,0.0390625,-0.0859375,-0.0625,-0.0078125,-0.0390625,-0.03125,0.1328125,-0.015625,-0.0390625,-0.046875,0.03125,0.0,0.0078125,-0.015625,-0.0078125,0.0078125,-0.0078125,-0.0,-0.0,-0.0078125,0.0234375,-0.046875,0.03125,0.09375,-0.078125,-0.0625,-0.046875,-0.0078125,-0.015625,-0.0234375,-0.078125,-0.078125,-0.0234375,0.03125,0.03125,0.03125,0.0078125,-0.015625,-0.0390625,-0.03125,-0.0859375,-0.078125,0.0546875,0.0390625,-0.0546875,0.0625,-0.046875,0.0078125,-0.015625,-0.0078125,-0.0546875,-0.0625,-0.015625,0.0546875,-0.046875,-0.0078125,0.015625,-0.0078125,-0.0078125,-0.015625,0.0,-0.0625,0.0234375,-0.0390625,-0.0234375,0.0234375,-0.0390625,-0.0078125,0.03125,-0.015625,0.0,-0.0703125,-0.046875,0.0078125,-0.0390625,0.0078125,0.0078125,0.0078125,-0.03125,-0.0234375,-0.015625,0.03125,-0.015625,-0.0234375,-0.0234375,0.0546875,0.0390625,-0.015625,0.046875,-0.0234375,-0.03125,-0.015625,-0.0546875,-0.046875,-0.0234375,0.015625,-0.03125,0.0234375,-0.0078125,0.0,0.0390625,0.0234375,-0.0625,-0.046875,-0.0234375,-0.046875,-0.03125,0.0625,0.0078125,0.1015625,0.0078125,0.0,0.0078125,-0.015625,-0.0078125,0.0078125,-0.0078125,-0.015625,-0.0078125,0.140625,0.109375,-0.015625,-0.0859375,-0.0703125,-0.0703125,-0.0390625,0.0078125,0.0078125,-0.03125,-0.015625,-0.046875,0.0234375,-0.03125,0.0859375,0.03125,-0.0078125,0.0078125,-0.0546875,-0.0859375,-0.03125,0.0078125,0.046875,0.015625,0.0234375,-0.015625,-0.0234375,0.03125,0.0234375,-0.0546875,-0.0390625,-0.0546875,0.0390625,-0.0234375,-0.0625,0.0234375,-0.0390625,0.0078125,-0.046875,0.0234375,-0.0,0.0390625,0.046875,0.0234375,-0.0,0.0546875,0.0390625,-0.0234375,-0.0078125,-0.0234375,0.03125,-0.0078125,-0.0078125,-0.03125,-0.03125,0.015625,-0.0234375,-0.0703125,-0.09375,0.1015625,-0.015625,-0.0625,0.046875,0.0390625,-0.0,-0.0234375,0.046875,-0.0546875,-0.0234375,-0.0625,-0.0390625,-0.0234375,0.015625,0.0625,0.0625,0.078125,0.046875,0.0703125,-0.03125,-0.09375,0.0234375,-0.0859375,0.0078125,-0.0234375,0.078125,0.0859375,0.0,0.0390625,0.0703125,0.0078125,0.015625,0.0859375,0.0390625,0.1171875,-0.0703125,-0.0390625,-0.03125,-0.078125,0.0,0.015625,-0.0625,0.0234375,0.0234375,-0.0,0.0625,0.0625,-0.0078125,-0.0078125,0.046875,-0.046875,0.03125,0.015625,-0.0,0.0,0.03125,0.015625,0.03125,0.078125,-0.078125,0.015625,0.015625,-0.015625,0.0078125,-0.0390625,0.0234375,-0.03125,0.0390625,-0.03125,-0.015625,-0.0390625,-0.09375,-0.0,0.0234375,0.015625,0.015625,0.0390625,-0.0546875,-0.015625,-0.0,-0.0078125,-0.0234375,-0.0,-0.0390625,0.0390625,0.0078125,-0.0078125,0.0078125,-0.0078125,-0.015625,0.015625,-0.015625,0.015625,-0.0,0.015625,0.046875,-0.0078125,0.03125,-0.078125,-0.078125,-0.0390625,0.015625,0.125,0.03125,0.0234375,0.0234375,-0.0078125,-0.0234375,0.0,-0.0625,0.015625,0.0078125,-0.03125,-0.0078125,-0.0390625,0.015625,-0.0234375,-0.046875,0.0390625,-0.0,0.0234375,-0.0,0.0078125,-0.0078125,-0.0078125,-0.0078125,0.0,-0.0078125,-0.0078125,0.0078125,-0.0078125,-0.046875,-0.0234375,-0.0390625,-0.0234375,-0.015625,-0.0546875,0.109375,-0.0625,0.0,0.0234375,-0.015625,-0.0078125,-0.015625,0.03125,-0.0078125,0.046875,0.09375,0.0390625,-0.03125,-0.03125,0.0,-0.0234375,-0.0390625,-0.015625,-0.0625,0.0546875,0.015625,-0.03125,-0.0078125,0.0,-0.015625,-0.015625,-0.0234375,0.0078125,0.0390625,0.0625,-0.0390625,-0.0546875,0.0078125,0.0546875,-0.0078125,0.0546875,0.015625,-0.0625,-0.015625,-0.015625,0.0,-0.046875,-0.03125,0.0625,0.015625,0.0390625,0.0546875,0.0078125,0.0,0.0078125,-0.0234375,-0.0078125,0.015625,-0.0078125,-0.0078125,0.015625,-0.0,-0.0,-0.015625,-0.046875,-0.0390625,0.0,0.03125,-0.0390625,-0.0390625,-0.0234375,-0.0,0.0,-0.0078125,0.0078125,-0.0703125,-0.0078125,0.0546875,-0.0078125,-0.015625,-0.0,-0.0390625,0.03125,0.03125,0.0078125,0.0234375,-0.03125,-0.09375,-0.0078125,0.0078125,-0.0,0.0078125,-0.0078125,-0.0234375,-0.0078125,-0.0234375,-0.0078125,0.03125,0.0,0.0078125,-0.015625,0.015625,-0.0234375,-0.03125,0.0390625,0.03125,-0.015625,-0.0234375,0.0234375,-0.03125,-0.0078125,0.0078125,-0.0078125,0.03125,0.03125,-0.0390625,0.0234375,0.015625,0.0,-0.0703125,-0.0234375,-0.0078125,-0.0078125,0.0859375,-0.0234375,0.0078125,-0.0078125,-0.0625,-0.046875,0.0390625,0.0,0.0234375,-0.046875,-0.0078125,0.0078125,0.0234375,0.0,-0.0390625,0.0234375,0.03125,-0.0234375,0.015625,-0.015625,0.03125,-0.03125,0.015625,-0.0703125,-0.0390625,0.0390625,-0.0234375,0.0390625,-0.0546875,0.0234375,0.0546875,-0.015625,-0.015625,0.0,0.0078125,-0.0234375,-0.046875,-0.0546875,0.0078125,0.03125,-0.0546875,0.0078125,0.015625,0.0234375,-0.0234375,0.0859375,-0.015625,0.046875,0.0390625,-0.0078125,-0.078125,-0.1015625,0.1171875,-0.0390625,-0.0234375,0.0078125,-0.0234375,-0.03125,0.0,0.0078125,0.03125,0.015625,-0.03125,0.0390625,0.0390625,-0.03125,-0.0546875,0.046875,-0.0234375,-0.0234375,-0.03125,-0.0546875,-0.09375,0.0390625,-0.0234375,-0.0078125,-0.0625,0.015625,-0.0078125,-0.0234375,-0.046875,0.015625,-0.015625,0.046875,-0.0078125,-0.0,-0.0078125,0.015625,0.015625,0.0078125,-0.046875,-0.0078125,0.0234375,-0.0234375,-0.0390625,-0.0234375,0.015625,0.03125,0.0390625,0.03125,-0.015625,0.0078125,0.0078125,-0.03125,0.03125,-0.0,-0.046875,-0.0390625,0.0234375,-0.0,0.0390625,0.0078125,0.0,0.015625,-0.0625,-0.0234375,0.078125,-0.0078125,-0.0078125,0.0,0.015625,-0.015625,-0.015625,0.015625,-0.0078125,-0.0,0.0078125,0.015625,-0.0234375,-0.0234375,-0.046875,-0.015625,-0.03125,0.0,0.015625,0.03125,0.0,0.0234375,-0.0,-0.03125,-0.0859375,0.0078125,-0.0078125,-0.0,0.015625,0.03125,-0.0078125,0.03125,-0.03125,-0.078125,-0.0625,0.0390625,0.015625,0.015625,0.0078125,0.015625,-0.0,-0.0078125,-0.0078125,-0.0078125,0.0078125,-0.0078125,-0.0,0.03125,-0.046875,0.078125,-0.0546875,-0.078125,-0.0,-0.046875,-0.1015625,0.0078125,-0.015625,-0.0625,-0.015625,0.0078125,0.03125,-0.046875,0.078125,0.09375,-0.046875,-0.015625,0.046875,0.2421875,-0.0390625,-0.0546875,-0.046875,-0.0390625,-0.0859375,-0.0234375,-0.0390625,-0.0546875,-0.0390625,-0.0234375,-0.0234375,-0.03125,-0.0234375,0.0234375,-0.0,-0.0390625,0.0078125,-0.0078125,0.0,-0.0625,-0.0078125,0.0390625,-0.0078125,0.0234375,-0.0234375,-0.015625,0.0234375,0.0390625,0.09375,0.0703125,-0.0234375,-0.0078125,-0.0546875,0.0,0.0546875,0.0,0.0,0.046875,0.03125,-0.0078125,-0.0078125,-0.0078125,0.0390625,-0.0078125,-0.0078125,-0.0625,-0.046875,0.015625,0.0,-0.0078125,-0.015625,-0.0390625,0.0703125,0.0234375,-0.0390625,-0.0625,0.0234375,0.0390625,0.0390625,0.015625,-0.015625,-0.015625,0.078125,0.015625,-0.0625,-0.0703125,0.03125,0.03125,0.046875,-0.0,-0.0234375,-0.0078125,0.015625,0.0078125,-0.0,0.0078125,0.0390625,-0.0,0.0078125,-0.0078125,-0.0078125,-0.046875,0.046875,-0.0,0.0,-0.0234375,-0.0078125,0.015625,-0.015625,-0.0078125,-0.0078125,0.109375,0.0390625,-0.046875,-0.0625,-0.046875,0.03125,-0.03125,0.015625,-0.015625,-0.0078125,0.0703125,-0.03125,-0.0078125,0.0078125,-0.0,-0.0390625,-0.03125,0.0078125,0.015625,-0.0078125,0.0390625,0.015625,0.046875,0.0234375,-0.0234375,-0.0234375,0.0625,-0.015625,-0.03125,0.0,-0.0078125,0.015625,-0.0234375,0.0234375,-0.0,-0.0390625,-0.0234375,0.1171875,-0.0078125,-0.03125,0.078125,0.0390625,-0.109375,0.1484375,-0.046875,-0.0546875,0.0234375,-0.1015625,-0.0390625,-0.0234375,-0.0,-0.0234375,0.0,0.0,-0.0546875,0.078125,-0.0078125,-0.0625,0.0078125,-0.015625,-0.0,0.015625,0.0078125,-0.046875,0.109375,-0.0078125,-0.0,-0.0546875,-0.0390625,-0.0234375,-0.03125,0.046875,0.0703125,0.015625,-0.03125,0.015625,-0.0625,-0.09375,-0.0234375,-0.03125,0.0,-0.109375,0.078125,0.0859375,-0.0390625,0.0234375,-0.0078125,0.0546875,0.015625,-0.0234375,-0.125,-0.0234375,0.03125,-0.0078125,-0.0703125,-0.0078125,0.0703125,-0.0,0.0078125,-0.1015625,0.0234375,-0.0234375,-0.03125,0.0234375,0.0390625,-0.0390625,0.046875,-0.0546875,0.0390625,0.03125,-0.046875,0.0078125,-0.0078125,0.0390625,0.0078125,0.015625,0.078125,-0.046875,0.015625,-0.0078125,-0.03125,0.0078125,-0.015625,0.0390625,-0.0,-0.0390625,0.1171875,-0.0,-0.046875,0.0390625,0.0234375,0.0078125,0.0,0.0078125,0.0078125,0.015625,0.0,0.015625,0.0078125,-0.0,0.0390625,0.046875,-0.046875,0.046875,-0.0234375,-0.0703125,-0.03125,-0.0703125,0.03125,0.0078125,-0.0078125,0.0390625,-0.0390625,-0.046875,-0.0234375,-0.0390625,-0.0234375,-0.0390625,0.0234375,-0.015625,-0.0234375,-0.0078125,-0.03125,-0.03125,0.046875,0.0078125,-0.0234375,-0.0078125,0.0078125,0.0078125,-0.0078125,-0.0,-0.0,0.0078125,-0.015625,-0.0078125,-0.0390625,0.046875,-0.046875,-0.015625,0.0703125,-0.015625,-0.0234375,-0.03125,0.0625,0.0859375,-0.0390625,0.015625,-0.0625,-0.0234375,-0.0078125,-0.0078125,0.0859375,0.0546875,-0.015625,-0.0703125,0.0078125,-0.078125,-0.0546875,-0.0703125,0.109375,0.0625,-0.0390625,-0.015625,-0.0,-0.0234375,0.015625,-0.03125,0.0,-0.03125,-0.015625,0.0234375,0.0234375,-0.0234375,-0.046875,-0.015625,0.0625,-0.0625,0.0078125,0.0390625,-0.0078125,-0.03125,-0.0234375,-0.0234375,0.0234375,-0.0234375,0.0,0.0234375,-0.015625,-0.0,-0.0,-0.015625,0.0078125,0.03125,-0.0234375,0.015625,-0.0078125,0.03125,0.03125,0.0,-0.0390625,-0.0,-0.03125,-0.0546875,0.0390625,0.0234375,-0.0078125,-0.03125,0.0234375,-0.0625,0.0234375,0.03125,0.0703125,-0.03125,-0.0234375,0.046875,-0.0078125,0.0234375,0.0,-0.0,0.0625,0.0390625,0.0390625,-0.015625,-0.078125,0.015625,-0.0078125,-0.015625,-0.0078125,-0.0078125,0.015625,0.0078125,0.0,0.0390625,0.0078125,-0.0078125,-0.015625,-0.0078125,-0.015625,-0.0234375,-0.0078125,-0.0,-0.03125,0.0078125,-0.03125,-0.0234375,0.0078125,0.0390625,-0.0234375,-0.03125,0.0234375,0.015625,-0.0546875,-0.015625,0.0,-0.0390625,-0.0390625,-0.0625,-0.015625,-0.0078125,0.03125,0.03125,-0.015625,-0.0859375,0.015625,-0.046875,0.03125,0.0625,0.0078125,0.1328125,-0.0390625,0.015625,0.015625,-0.0078125,0.0625,-0.0234375,0.0078125,-0.0625,0.0390625,0.015625,0.0078125,0.0546875,-0.0078125,0.0546875,-0.109375,-0.0234375,-0.0234375,-0.0234375,-0.0078125,-0.0390625,-0.0234375,-0.0390625,-0.03125,0.0234375,0.0546875,-0.0,-0.0625,-0.0390625,-0.0078125,-0.015625,-0.0078125,0.0234375,-0.015625,-0.0546875,0.03125,0.0234375,-0.0703125,0.078125,-0.0234375,-0.0234375,-0.03125,-0.0625,0.0,0.03125,-0.015625,-0.0546875,-0.0234375,-0.015625,-0.0078125,0.015625,-0.046875,0.0078125,-0.0,-0.015625,0.0546875,-0.015625,-0.0234375,-0.0390625,0.0390625,0.0234375,0.03125,-0.03125,0.0078125,-0.09375,0.03125,-0.0546875,0.0078125,-0.0078125,-0.1015625,0.0390625,-0.09375,0.09375,0.0078125,0.0546875,0.0078125,0.0078125,-0.0078125,-0.03125,0.0234375,-0.0078125,-0.0625,0.0234375,-0.0078125,0.0390625,0.015625,0.046875,0.0,-0.0,-0.0,-0.0234375,0.0390625,-0.0546875,0.03125,-0.015625,-0.046875,0.0234375,0.0703125,-0.0234375,0.0078125,-0.0625,-0.015625,0.0703125,0.0078125,-0.0546875,0.03125,-0.015625,-0.015625,-0.0234375,-0.0,-0.015625,-0.015625,-0.0,-0.0078125,0.0078125,-0.0,-0.0078125,0.0078125,-0.0,0.03125,-0.0546875,0.015625,0.1015625,0.015625,-0.03125,0.0234375,-0.078125,0.0078125,-0.046875,-0.0625,0.0546875,0.03125,0.0546875,-0.015625,0.046875,0.0625,0.015625,0.0078125,0.015625,0.015625,-0.0546875,0.046875,-0.0234375,0.03125,0.0,-0.0078125,0.0,-0.0,-0.015625,-0.0078125,-0.0078125,0.0,0.0078125,0.0078125,-0.0078125,-0.0390625,0.0859375,0.0,-0.0546875,-0.0,0.0234375,0.0078125,-0.046875,-0.0390625,-0.046875,-0.0859375,0.0078125,-0.046875,-0.0390625,-0.0234375,-0.0546875,-0.0,0.015625,0.0078125,-0.0078125,-0.046875,0.03125,0.015625,-0.0625,-0.03125,0.046875,0.03125,0.0078125,0.015625,0.0234375,-0.0078125,0.015625,0.046875,-0.015625,-0.015625,-0.03125,0.0390625,0.0390625,0.03125,-0.03125,-0.0625,-0.0,-0.0,-0.0625,0.0,-0.0390625,-0.0703125,0.03125,-0.0,-0.015625,0.0078125,0.0078125,-0.0234375,-0.0078125,-0.0234375,0.0078125,0.0,-0.015625,0.0,0.0078125,-0.015625,0.03125,-0.0078125,0.0078125,0.03125,0.03125,-0.0078125,-0.0078125,0.0390625,-0.0078125,-0.015625,0.0078125,0.0,0.0625,-0.0078125,-0.0546875,-0.0390625,-0.015625,0.0703125,0.0078125,0.0078125,-0.0625,0.0859375,-0.0703125,-0.03125,0.03125,0.0234375,0.0625,-0.0546875,-0.015625,-0.0234375,-0.0,-0.0,0.0078125,0.0,0.03125,-0.015625,-0.015625,0.0,0.0078125,-0.0546875,0.0078125,0.0703125,-0.015625,-0.015625,-0.0390625,0.015625,0.0,-0.0,0.015625,-0.0078125,-0.046875,-0.0234375,-0.0078125,-0.0078125,0.0234375,-0.03125,0.1484375,0.015625,-0.0546875,-0.078125,0.0078125,-0.0546875,-0.046875,-0.03125,0.0,-0.0078125,-0.0234375,-0.046875,-0.0234375,0.09375,0.015625,0.0078125,0.0078125,-0.0234375,0.03125,-0.078125,-0.0546875,0.0546875,0.078125,-0.0,-0.078125,-0.015625,-0.046875,-0.0234375,-0.015625,-0.0078125,-0.03125,-0.0390625,-0.0546875,0.015625,-0.0390625,0.0234375,-0.046875,-0.0390625,-0.03125,0.015625,0.0625,0.0390625,-0.0390625,-0.015625,0.0234375,0.015625,0.0390625,-0.0390625,0.0,0.0234375,0.0234375,0.0,-0.015625,0.015625,-0.046875,-0.0,0.0390625,0.046875,0.015625,-0.0078125,-0.0625,0.0234375,0.0625,-0.015625,0.0390625,-0.03125,0.015625,-0.0,0.03125,-0.0703125,-0.046875,0.0078125,0.015625,0.109375,0.03125,0.015625,-0.0390625,-0.0234375,0.046875,-0.0234375,-0.0390625,0.0234375,0.1171875,0.0078125,-0.046875,-0.03125,-0.0625,0.03125,0.0078125,-0.0234375,-0.0234375,-0.0078125,0.0546875,0.0234375,-0.1015625,0.0234375,-0.0234375,0.0078125,-0.0078125,-0.0625,-0.0234375,-0.0546875,0.0078125,-0.015625,-0.03125,0.0546875,-0.0,-0.0,-0.0078125,-0.0703125,-0.0,0.03125,0.0,-0.0234375,-0.0234375,0.0,-0.0,-0.015625,-0.046875,0.015625,-0.015625,0.03125,-0.0234375,-0.03125,-0.0078125,0.046875,0.0,0.0078125,-0.0078125,0.0,0.0234375,0.0078125,-0.0,0.0234375,-0.015625,-0.0234375,-0.0078125,-0.0546875,-0.0078125,-0.0078125,-0.0234375,-0.0234375,-0.0390625,0.015625,-0.0078125,0.0546875,0.0,-0.0078125,0.046875,-0.0390625,-0.015625,0.03125,0.03125,-0.0078125,0.0234375,0.0234375,-0.0078125,-0.015625,-0.0859375,-0.0390625,-0.0625,0.0234375,0.0078125,-0.0078125,0.0078125,0.0,0.0078125,0.0078125,-0.0078125,0.0078125,-0.0,-0.0078125,-0.015625,-0.0078125,-0.0234375,-0.015625,0.0390625,-0.046875,0.0546875,-0.0,-0.0078125,0.0078125,-0.015625,-0.015625,0.015625,-0.1015625,-0.015625,0.0859375,0.0234375,0.0078125,-0.0,0.03125,-0.0078125,0.0,-0.0390625,-0.015625,-0.0078125,0.0703125,-0.0078125,-0.015625,0.0234375,0.0078125,0.0078125,0.0546875,0.015625,-0.046875,-0.0078125,-0.015625,0.015625,0.03125,-0.015625,-0.0078125,0.0078125,-0.015625,0.09375,0.0703125,-0.015625,-0.0234375,-0.0234375,-0.015625,0.0078125,0.03125,-0.0078125,0.0390625,0.0234375,0.0078125,-0.015625,0.0078125,-0.015625,-0.015625,-0.03125,-0.015625,0.015625,-0.0078125,-0.0078125,-0.0,-0.0234375,-0.0234375,-0.0078125,-0.03125,-0.0,-0.0,0.0390625,-0.0078125,0.015625,0.0234375,-0.015625,0.0,-0.046875,-0.015625,0.03125,-0.0234375,-0.015625,-0.046875,0.0625,-0.03125,-0.046875,-0.015625,-0.015625,-0.0703125,-0.0546875,0.0078125,-0.0078125,-0.0,0.0078125,0.0078125,-0.0,-0.015625,-0.0078125,-0.015625,0.0,0.015625,-0.0234375,-0.015625,0.0078125,0.0390625,0.0078125,0.03125,0.0546875,-0.015625,0.0546875,0.0078125,-0.015625,0.0234375,0.03125,-0.0078125,0.0703125,-0.0234375,-0.015625,-0.0078125,0.0,-0.0,-0.0078125,-0.109375,-0.0,0.0078125,0.046875,-0.015625,0.0234375,0.0078125,-0.0234375,-0.0234375,-0.046875,-0.0078125,0.0078125,-0.015625,-0.015625,-0.0546875,0.03125,-0.0078125,-0.078125,-0.0390625,-0.015625,-0.046875,-0.0390625,-0.0078125,0.0,0.0078125,-0.03125,-0.0234375,0.0390625,-0.0390625,0.0078125,-0.0078125,-0.0234375,0.0234375,0.0390625,-0.0,0.0546875,-0.03125,-0.0078125,0.0390625,0.03125,-0.0078125,-0.015625,0.0390625,-0.015625,-0.015625,0.0703125,0.015625,0.0625,-0.03125,0.0078125,-0.0078125,0.015625,-0.015625,-0.015625,-0.0234375,-0.0078125,0.015625,-0.046875,-0.0078125,-0.0234375,-0.0078125,-0.0078125,-0.0234375,-0.03125,-0.0234375,-0.0234375,0.0234375,-0.0234375,-0.015625,0.0390625,-0.046875,-0.0078125,-0.015625,-0.015625,-0.015625,-0.015625,-0.0,0.0390625,0.0390625,-0.015625,0.0078125,-0.0390625,-0.015625,-0.0390625,0.0078125,-0.015625,-0.03125,-0.015625,-0.03125,-0.0625,-0.03125,-0.03125,-0.015625,0.015625,-0.0078125,0.0078125,0.046875,-0.015625,-0.0703125,-0.0546875,-0.03125,0.0234375,-0.0546875,-0.03125,0.046875,-0.03125,-0.0234375,0.0,-0.0234375,-0.0078125,0.046875,-0.0078125,0.0546875,0.046875,0.046875,-0.015625,-0.046875,0.0078125,0.0390625,0.0078125,-0.0390625,-0.0078125,-0.0078125,0.0,-0.0,0.0078125,0.0078125,-0.0078125,0.015625,0.0,-0.0625,-0.015625,-0.0234375,0.0703125,-0.0234375,-0.0078125,-0.0234375,-0.03125,0.0234375,0.0,0.0,-0.0234375,0.0078125,-0.0546875,0.03125,-0.015625,-0.046875,0.03125,-0.015625,0.03125,-0.046875,0.0078125,-0.015625,-0.015625,-0.0078125,0.03125,-0.0234375,-0.0078125,-0.015625,-0.0078125,0.0,0.0078125,0.0,-0.0078125,0.0,-0.0078125,-0.0625,-0.015625,0.0,-0.0390625,-0.09375,-0.0078125,0.09375,0.015625,-0.0390625,0.109375,-0.046875,-0.0390625,-0.0078125,-0.0703125,-0.046875,0.015625,0.0078125,-0.046875,0.0078125,0.0703125,-0.0078125,-0.0546875,-0.0546875,-0.046875,0.0390625,0.03125,0.0390625,0.0078125,-0.0390625,-0.0234375,0.0078125,0.015625,-0.03125,0.0625,0.0078125,0.015625,0.0078125,0.046875,0.03125,-0.1171875,-0.0546875,-0.03125,0.0234375,0.0234375,-0.0078125,-0.0234375,-0.046875,-0.0234375,0.0234375,0.0546875,-0.015625,-0.015625,-0.0,-0.0390625,0.0546875,0.015625,-0.0234375,-0.03125,-0.0078125,-0.0078125,-0.0078125,0.015625,-0.0,-0.0078125,-0.0234375,0.0078125,-0.0234375,0.0234375,0.015625,0.0390625,-0.0078125,0.0078125,-0.0234375,-0.0390625,-0.0078125,-0.046875,-0.015625,-0.078125,0.0703125,0.0625,-0.046875,-0.0234375,0.0390625,-0.0625,-0.0,-0.0546875,-0.046875,0.0078125,0.109375,-0.0,-0.0078125,-0.0,0.0,0.015625,0.0078125,0.0,-0.015625,0.015625,0.0,0.0234375,-0.0625,-0.015625,0.0546875,0.015625,-0.0078125,-0.0390625,-0.015625,-0.0078125,0.0078125,-0.0078125,0.015625,-0.015625,-0.046875,0.03125,-0.0078125,-0.03125,0.0234375,0.0,-0.0390625,-0.0078125,0.140625,0.0703125,0.0078125,0.046875,0.0859375,-0.0703125,-0.09375,0.0234375,0.046875,0.0625,-0.0859375,0.0234375,0.140625,0.03125,0.015625,0.0546875,-0.0078125,-0.015625,-0.0546875,0.0390625,-0.03125,-0.0546875,0.0859375,-0.0390625,0.03125,0.03125,0.046875,-0.0703125,0.046875,-0.0234375,-0.046875,0.015625,-0.0,-0.0390625,-0.015625,-0.0078125,0.125,0.0078125,0.015625,-0.1640625,-0.0078125,-0.0,0.0546875,-0.0078125,0.0234375,-0.015625,0.0390625,-0.015625,-0.0,-0.0390625,0.0,0.0078125,0.0234375,0.015625,-0.0625,-0.015625,0.0078125,-0.046875,-0.0546875,-0.0234375,0.0390625,-0.0625,-0.0234375,0.0,-0.03125,-0.0234375,0.1015625,0.03125,0.0,-0.0546875,-0.09375,-0.015625,0.0078125,-0.0234375,-0.03125,0.0546875,-0.015625,-0.03125,-0.0625,-0.0390625,0.015625,0.0625,-0.0390625,0.0078125,-0.078125,-0.0234375,-0.0390625,-0.0546875,-0.046875,-0.03125,0.0078125,-0.0234375,-0.0546875,-0.046875,0.015625,-0.015625,-0.015625,0.03125,0.015625,0.0546875,0.0390625,-0.03125,0.015625,0.0078125,-0.03125,0.0390625,-0.046875,0.0078125,0.0078125,-0.0,-0.0078125,-0.015625,0.0234375,-0.0078125,-0.03125,-0.0078125,-0.0390625,0.0078125,0.0625,0.0234375,-0.0078125,-0.03125,-0.0390625,0.015625,0.0078125,-0.0,0.0078125,-0.015625,0.0078125,-0.015625,-0.0078125,0.0078125,-0.0390625,-0.015625,0.0546875,0.015625,0.015625,0.0,0.0,0.0078125,0.015625,0.0078125,0.0078125,0.0234375,0.015625,0.0078125,-0.046875,0.0,0.0234375,-0.0,-0.0078125,-0.015625,0.0703125,-0.0,-0.046875,-0.015625,-0.0,-0.03125,0.0078125,0.0078125,0.0,0.015625,0.0078125,-0.0078125,-0.0078125,0.0,-0.0,-0.0078125,0.0234375,-0.015625,-0.03125,-0.0703125,-0.046875,-0.046875,-0.0,0.0,-0.0078125,0.03125,0.0234375,0.015625,-0.0234375,-0.0859375,0.0625,-0.015625,-0.015625,-0.0234375,0.0859375,0.078125,0.0546875,-0.0234375,-0.03125,-0.0390625,-0.015625,0.015625,0.0234375,-0.0078125,-0.015625,-0.0078125,-0.015625,-0.03125,-0.015625,-0.015625,-0.015625,-0.015625,-0.03125,0.0546875,-0.0234375,-0.015625,0.0234375,0.0546875,-0.0078125,-0.015625,0.0,0.0390625,0.0,0.0234375,-0.0234375,-0.0859375,0.0078125,-0.015625,-0.015625,-0.0078125,0.0078125,0.0,0.0078125,0.015625,0.0078125,-0.0234375,0.015625,-0.0078125,-0.0078125,-0.0078125,0.015625,0.0390625,-0.0078125,-0.0390625,0.0625,0.0,0.0078125,0.0234375,-0.015625,0.03125,-0.015625,0.0078125,0.0234375,0.0078125,-0.0078125,-0.015625,-0.0,0.015625,-0.078125,0.078125,-0.046875,-0.0234375,-0.03125,-0.03125,-0.0234375,-0.0234375,-0.015625,-0.0234375,0.015625,-0.0078125,-0.0078125,0.015625,0.0078125,-0.0078125,0.0,0.015625,0.0,-0.015625,-0.0078125,-0.0390625,-0.015625,0.015625,-0.03125,-0.015625,-0.03125,-0.0234375,-0.0625,0.0,0.0078125,0.0,0.0078125,-0.015625,0.015625,0.0390625,0.0546875,0.0234375,-0.0,-0.0546875,0.03125,-0.015625,-0.0546875,-0.0546875,0.0,0.0,-0.046875,-0.0546875,0.0234375,0.046875,-0.0,-0.0,0.0390625,-0.015625,-0.03125,-0.015625,0.0078125,-0.09375,-0.03125,-0.015625,-0.078125,-0.0390625,-0.015625,0.0625,0.046875,0.0234375,0.015625,-0.015625,-0.0,-0.0234375,0.0,0.0078125,-0.1015625,0.1171875,0.0859375,-0.0390625,-0.0234375,-0.015625,-0.0390625,-0.015625,-0.03125,-0.0390625,-0.0234375,-0.0234375,-0.09375,0.03125,-0.0,-0.015625,-0.0390625,0.046875,0.0,0.0625,0.0234375,-0.09375,0.0546875,-0.0078125,-0.015625,-0.0078125,-0.0234375,-0.0234375,-0.03125,0.0390625,-0.0234375,0.015625,0.015625,0.015625,0.0078125,-0.0078125,-0.0703125,-0.015625,0.0,0.0,-0.0234375,-0.0078125,0.015625,-0.0234375,-0.0234375,-0.1015625,-0.0625,0.0234375,0.0859375,0.0625,-0.015625,-0.03125,-0.0078125,-0.0390625,0.0625,-0.0234375,-0.0703125,0.0390625,-0.0390625,0.0078125,-0.0390625,-0.0234375,0.0,-0.0859375,-0.0,0.0234375,0.015625,0.0703125,-0.015625,0.0234375,0.0546875,-0.046875,0.046875,-0.03125,-0.03125,0.0078125,-0.0078125,-0.0078125,-0.0078125,-0.015625,-0.0078125,-0.0078125,-0.0,0.0390625,0.09375,0.0,-0.0390625,-0.015625,-0.0234375,-0.0,-0.015625,-0.0078125,-0.0,-0.0234375,0.0,-0.0078125,0.0078125,-0.0078125,-0.015625,0.0078125,-0.0390625,-0.0078125,0.046875,0.015625,0.03125,-0.015625,0.0234375,-0.03125,-0.015625,-0.03125,-0.0,-0.015625,-0.0703125,0.046875,0.0078125,0.109375,0.015625,-0.0390625,0.015625,-0.0546875,-0.0625,-0.0703125,0.0234375,-0.0703125,0.046875,0.0078125,0.0,-0.0078125,0.0078125,-0.0078125,0.0078125,-0.0,-0.0078125,0.0078125,-0.046875,0.0234375,-0.0625,-0.046875,-0.015625,0.03125,-0.046875,0.0078125,0.078125,-0.015625,-0.0390625,0.0,-0.0390625,-0.0390625,0.03125,0.0,0.0078125,-0.0,-0.0,-0.0546875,-0.0390625,-0.03125,0.203125,-0.0078125,-0.0859375,0.03125,-0.0625,-0.0234375,-0.0078125,-0.046875,-0.0703125,0.09375,-0.0390625,0.0,-0.0,0.0,0.0546875,-0.0390625,-0.0234375,0.0234375,-0.0546875,-0.0078125,-0.015625,-0.0390625,-0.0234375,0.0078125,-0.0234375,-0.03125,-0.0,-0.046875,-0.0078125,-0.0234375,-0.0625,-0.03125,0.015625,0.015625,-0.015625,0.015625,0.0078125,-0.0234375,-0.0078125,0.03125,-0.0234375,-0.0078125,-0.0234375,-0.0078125,-0.015625,-0.0390625,-0.046875,0.015625,-0.125,0.015625,0.0390625,-0.0,0.0078125,-0.0546875,-0.0703125,-0.0234375,0.0390625,0.0703125,0.0078125,0.03125,0.0078125,0.0078125,0.0078125,0.046875,0.015625,-0.0234375,0.015625,0.0234375,-0.0078125,-0.0078125,-0.0,0.015625,0.0078125,-0.0078125,-0.0078125,0.03125,-0.0078125,-0.0234375,0.0,-0.015625,-0.0546875,0.0625,-0.015625,-0.015625,0.0703125,-0.0,-0.0859375,-0.015625,-0.078125,0.1015625,-0.046875,0.09375,0.0546875,0.046875,0.0,0.015625,-0.0390625,0.03125,-0.015625,-0.046875,0.015625,-0.0234375,-0.078125,-0.0703125,-0.015625,-0.0078125,-0.0546875,-0.0390625,-0.0390625,0.015625,0.03125,-0.078125,-0.015625,0.015625,-0.0078125,-0.015625,-0.046875,-0.046875,-0.03125,-0.0625,-0.0,-0.0234375,0.015625,0.0078125,0.015625,0.0234375,-0.03125,0.0078125,0.0234375,0.046875,-0.03125,-0.015625,-0.0625,-0.046875,0.0234375,-0.1640625,0.09375,0.078125,-0.1171875,0.0390625,-0.0078125,-0.0078125,-0.0078125,-0.015625,0.0703125,-0.0078125,0.0234375,0.0625,-0.0390625,0.03125,0.03125,0.046875,-0.1171875,-0.09375,-0.03125,0.0546875,0.0078125,0.015625,-0.0078125,-0.0234375,-0.0390625,0.078125,-0.109375,-0.046875,0.0078125,0.0078125,0.0,-0.015625,-0.0234375,-0.0859375,-0.0,0.015625,-0.0078125,0.09375,-0.015625,0.0390625,0.0390625,0.0078125,0.0234375,-0.046875,-0.1640625,-0.046875,-0.0,-0.015625,0.0234375,-0.015625,-0.0234375,-0.015625,-0.0234375,-0.1484375,-0.03125,0.015625,-0.015625,0.0546875,0.0078125,0.0078125,0.0390625,0.0546875,-0.1328125,0.03125,0.0,0.1328125,0.015625,-0.015625,-0.0703125,0.0078125,0.046875,-0.0625,0.078125,-0.078125,-0.0390625,0.0078125,-0.0625,0.046875,0.09375,-0.0078125,-0.0234375,-0.0625,0.0078125,0.0078125,-0.0625,0.0078125,0.015625,-0.0,-0.0078125,0.0234375,0.0078125,0.0,-0.015625,-0.015625,-0.015625,-0.0,-0.046875,0.0078125,0.046875,0.03125,0.03125,0.0078125,-0.0390625,-0.0078125,-0.0078125,0.015625,0.0546875,-0.046875,0.046875,0.015625,-0.0859375,-0.0078125,0.0078125,-0.0390625,-0.046875,-0.0078125,0.1015625,0.0078125,-0.015625,-0.015625,-0.0078125,0.015625,0.0078125,0.03125,-0.0078125,-0.0,-0.0078125,0.0078125,0.0,-0.0078125,-0.0078125,-0.0625,-0.046875,-0.015625,0.1171875,-0.0546875,-0.0234375,0.0390625,0.03125,-0.03125,-0.0859375,0.15625,-0.046875,-0.03125,0.078125,-0.0390625,-0.1328125,-0.015625,0.015625,-0.0078125,-0.0234375,0.0390625,0.03125,0.015625,0.0078125,0.0078125,0.078125,0.0078125,0.015625,0.0703125,0.0,-0.0625,-0.03125,-0.0,0.03125,0.0,0.015625,-0.0,0.0078125,-0.03125,-0.015625,-0.0546875,-0.0078125,0.0078125,0.109375,-0.0234375,0.0625,0.0390625,-0.015625,0.0078125,-0.0234375,0.0234375,-0.015625,-0.0078125,0.015625,-0.0234375,0.015625,0.0,-0.0234375,-0.015625,-0.0078125,0.015625,-0.015625,0.0078125,-0.0234375,-0.046875,-0.046875,0.1171875,0.015625,-0.03125,-0.0078125,-0.0390625,-0.0078125,-0.0078125,-0.0859375,-0.0625,-0.0234375,0.125,-0.0078125,-0.0078125,-0.0078125,0.0,-0.0390625,0.09375,-0.0078125,0.0078125,0.03125,0.0078125,0.0234375,-0.046875,0.015625,0.0,-0.015625,-0.0,-0.0234375,-0.0,0.0,-0.015625,-0.015625,-0.0234375,-0.0234375,-0.0078125,0.0234375,-0.0234375,-0.03125,0.0234375,0.03125,-0.0078125,-0.0078125,-0.0078125,-0.0703125,-0.0078125,0.0078125,-0.0234375,-0.03125,0.0078125,-0.0390625,0.015625,0.046875,-0.0390625,-0.015625,-0.03125,0.078125,-0.0390625,0.078125,-0.046875,0.0078125,0.0390625,-0.0703125,-0.0390625,0.0546875,0.0546875,-0.03125,-0.0234375,0.03125,-0.0078125,0.03125,0.0234375,-0.015625,0.0234375,-0.078125,-0.0078125,-0.03125,0.0390625,-0.015625,0.0234375,-0.1015625,-0.0078125,-0.1015625,-0.0,0.0078125,0.0234375,-0.0859375,-0.0390625,0.0390625,-0.046875,-0.0234375,-0.0859375,0.0546875,-0.0,0.0390625,-0.0234375,-0.0078125,0.0625,0.0625,0.015625,0.03125,-0.0,0.0078125,-0.0,-0.03125,-0.0078125,0.0,-0.09375,0.015625,-0.03125,-0.0,0.015625,0.0234375,0.0546875,-0.0,0.03125,0.0703125,-0.03125,0.0078125,-0.046875,-0.0625,-0.0546875,0.0078125,0.0078125,-0.015625,0.046875,-0.0,0.0390625,0.03125,-0.0078125,-0.0390625,-0.0625,-0.0078125,-0.078125,-0.0625,-0.015625,-0.0234375,-0.015625,0.0,0.0546875,0.109375,-0.0234375,-0.015625,-0.0703125,-0.03125,-0.0234375,0.015625,-0.046875,-0.0078125,-0.0078125,0.0,0.078125,-0.0234375,-0.03125,0.015625,0.0390625,-0.0234375,-0.046875,-0.078125,-0.0625,0.0078125,0.171875,-0.046875,-0.1171875,-0.015625,0.0078125,-0.0078125,0.03125,-0.0546875,0.109375,0.1015625,0.03125,0.0859375,0.0078125,0.0078125,-0.0078125,-0.03125,0.015625,0.0078125,0.0,0.015625,-0.0078125,-0.0,0.0,0.0078125,0.0,0.0625,0.03125,0.046875,-0.03125,0.0078125,0.0078125,-0.0078125,-0.03125,-0.015625,0.0390625,0.0234375,-0.0625,0.0390625,0.0390625,-0.0625,0.015625,-0.015625,-0.0390625,-0.015625,-0.0234375,-0.0625,0.0234375,-0.046875,0.1015625,-0.0,0.0234375,-0.0234375,-0.015625,-0.0078125,-0.0078125,-0.0078125,0.0078125,0.0078125,0.015625,-0.015625,-0.0,0.109375,0.046875,-0.03125,-0.0078125,-0.046875,-0.015625,0.0078125,-0.046875,-0.0,0.03125,0.015625,0.0703125,-0.0546875,0.0,-0.0703125,-0.0234375,-0.0078125,-0.0078125,-0.03125,-0.046875,0.078125,-0.0703125,-0.015625,0.0234375,0.015625,-0.0234375,-0.015625,-0.0234375,0.0078125,0.0546875,0.0,-0.0234375,-0.0390625,-0.0078125,-0.03125,-0.0078125,-0.0390625,-0.0390625,0.1015625,-0.0078125,0.015625,-0.0,-0.0,0.03125,-0.03125,-0.0390625,0.015625,-0.0390625,-0.0,-0.0078125,-0.0234375,0.0078125,0.015625,0.015625,0.0234375,-0.03125,-0.0546875,0.015625,0.0,-0.0078125,0.0,0.0078125,-0.0078125,0.0546875,-0.0234375,-0.0390625,0.0234375,0.0078125,0.09375,-0.0,-0.015625,-0.015625,0.0,-0.0546875,0.0703125,-0.0625,0.0234375,0.0546875,-0.0234375,-0.015625,-0.0625,0.015625,0.0703125,-0.0078125,-0.046875,-0.0546875,-0.0234375,-0.015625,-0.015625,-0.0234375,-0.0078125,-0.0,0.015625,-0.015625,-0.015625,0.015625,-0.0,0.015625,0.015625,0.046875,-0.0625,-0.0,-0.0,0.0078125,-0.0078125,0.015625,-0.0390625,-0.0078125,-0.0234375,-0.0,-0.0859375,0.0625,0.0390625,-0.0546875,-0.0078125,-0.03125,-0.0078125,-0.046875,0.03125,0.0625,-0.078125,-0.046875,0.015625,-0.0234375,-0.0390625,-0.0234375,0.0234375,-0.109375,0.0703125,-0.0078125,0.0078125,0.0546875,-0.0390625,-0.03125,-0.015625,-0.0625,-0.0234375,0.0234375,0.0234375,-0.078125,-0.046875,-0.03125,-0.0546875,-0.0,0.0625,0.078125,0.0078125,-0.078125,0.0,0.03125,-0.0234375,-0.0390625,0.0078125,0.0390625,-0.046875,-0.0078125,-0.0234375,-0.0390625,-0.0859375,-0.0,-0.0546875,-0.0,-0.0390625,0.0078125,0.015625,-0.046875,0.0,0.0546875,-0.015625,-0.015625,-0.0,0.0078125,-0.0546875,-0.046875,-0.0703125,0.0390625,0.1171875,-0.015625,-0.015625,-0.015625,0.0234375,0.0234375,-0.015625,0.0390625,-0.046875,-0.0703125,-0.03125,-0.0234375,0.015625,-0.015625,0.109375,-0.0625,0.0859375,-0.0234375,-0.0234375,-0.0078125,-0.0234375,-0.015625,0.0859375,-0.1328125,-0.015625,0.078125,0.0390625,0.0234375,-0.0078125,0.03125,-0.0390625,0.0703125,0.046875,-0.0859375,0.0703125,-0.09375,0.0625,0.0078125,-0.0234375,-0.015625,0.046875,0.0234375,0.0625,0.0,-0.0703125,0.0078125,-0.0234375,0.0,-0.015625,0.0078125,-0.0,0.03125,0.0625,-0.0390625,-0.03125,-0.015625,-0.0390625,-0.0078125,-0.03125,0.109375,-0.046875,0.0234375,0.046875,0.0546875,-0.1171875,-0.015625,-0.0078125,-0.0078125,-0.0078125,-0.0,0.0,0.0,-0.015625,-0.0078125,-0.0078125,0.015625,0.0546875,0.0390625,0.0234375,-0.046875,-0.109375,-0.0546875,0.0078125,-0.0,-0.0234375,-0.03125,-0.03125,0.046875,-0.0078125,-0.03125,-0.0078125,-0.0234375,0.0390625,0.0703125,0.0234375,0.0078125,-0.0234375,-0.0,-0.1015625,-0.0390625,-0.0078125,0.0234375,-0.078125,0.0078125,0.015625,0.015625,-0.0,-0.0078125,-0.0078125,-0.0078125,-0.0078125,0.0,-0.0390625,-0.0703125,-0.0390625,0.0234375,-0.0859375,0.0625,-0.03125,0.03125,0.0546875,-0.03125,-0.0,-0.03125,-0.0,0.0234375,0.0078125,0.03125,0.0078125,0.0390625,0.0703125,0.03125,0.0078125,-0.078125,-0.0859375,-0.046875,0.03125,0.03125,-0.0234375,-0.0625,0.0390625,0.03125,-0.0234375,-0.046875,0.0625,-0.0234375,0.0703125,-0.0234375,0.0078125,-0.0078125,-0.0234375,-0.0625,0.0546875,-0.03125,0.015625,-0.109375,0.015625,0.0,-0.0078125,-0.03125,-0.015625,-0.03125,-0.0546875,-0.03125,0.0,-0.0078125,0.0234375,-0.0078125,-0.0078125,0.015625,0.0078125,0.0,-0.03125,0.0,0.03125,-0.015625,0.046875,0.0078125,-0.0625,-0.03125,-0.0390625,-0.015625,-0.0,-0.046875,-0.0703125,0.03125,-0.0859375,0.015625,-0.0703125,-0.03125,0.046875,-0.0,0.0078125,-0.0078125,0.015625,-0.0546875,0.0625,-0.0546875,-0.0,-0.03125,0.0390625,-0.109375,0.0,0.0078125,0.0078125,-0.0078125,-0.015625,0.0078125,0.015625,0.03125,0.015625,-0.015625,-0.015625,-0.015625,-0.046875,0.0,-0.0390625,-0.03125,0.0390625,0.0390625,0.03125,-0.03125,0.0625,0.0078125,-0.0234375,0.0234375,-0.046875,0.0390625,0.0390625,0.0,0.0234375,-0.0078125,0.0078125,-0.078125,-0.015625,0.0390625,0.015625,-0.03125,-0.0390625,0.09375,0.0078125,-0.125,-0.0078125,-0.1015625,-0.0078125,-0.078125,-0.0234375,-0.03125,-0.0390625,-0.0625,-0.0234375,-0.09375,0.015625,0.0625,0.1015625,0.015625,0.0390625,0.0234375,-0.0,0.0078125,-0.0390625,-0.0859375,0.0078125,-0.0390625,-0.015625,0.03125,-0.0234375,0.078125,-0.0234375,0.03125,-0.0078125,-0.046875,0.015625,-0.0390625,-0.0078125,0.0234375,-0.015625,-0.03125,-0.0078125,-0.0234375,0.015625,0.03125,0.0234375,-0.0,0.0625,0.03125,-0.078125,0.03125,-0.03125,-0.0546875,-0.0078125,0.0234375,-0.0078125,-0.046875,0.0546875,-0.0234375,-0.03125,-0.0390625,0.0234375,0.1171875,-0.0078125,0.15625,0.0078125,0.0234375,-0.0078125,0.078125,-0.03125,-0.078125,-0.0234375,-0.09375,0.015625,0.046875,-0.0390625,0.0625,0.046875,-0.0078125,-0.0078125,-0.09375,0.015625,0.03125,-0.0234375,0.0703125,-0.0546875,-0.015625,-0.0078125,0.078125,-0.0625,0.0703125,-0.0234375,0.0859375,-0.03125,-0.03125,0.046875,-0.0234375,-0.0234375,-0.015625,0.0078125,0.0859375,0.015625,0.046875,-0.015625,-0.0546875,0.015625,-0.0390625,0.015625,-0.0234375,0.125,0.0234375,0.0234375,-0.0234375,-0.1328125,-0.0078125,-0.03125,-0.0078125,-0.015625,0.0078125,0.03125,-0.0,0.0,-0.015625,-0.0078125,0.0078125,0.0078125,-0.0078125,0.0,-0.0546875,-0.0078125,-0.03125,0.015625,-0.046875,0.03125,0.015625,0.0625,0.0078125,0.0,0.0234375,0.0,-0.015625,-0.015625,0.0078125,0.0546875,0.0078125,-0.0234375,0.03125,-0.015625,0.015625,0.046875,0.0859375,-0.0078125,-0.0625,-0.0078125,0.0078125,0.0,-0.015625,-0.0078125,-0.015625,-0.0078125,-0.0078125,0.0078125,0.0078125,-0.0078125,-0.0546875,0.0078125,0.078125,-0.0390625,-0.078125,0.078125,-0.0234375,0.078125,0.0625,0.0703125,0.078125,-0.0390625,-0.078125,-0.1171875,-0.046875,-0.0390625,-0.0390625,0.0859375,-0.0078125,0.0234375,-0.046875,0.0390625,0.0234375,0.0,0.015625,-0.015625,-0.0390625,0.0078125,0.015625,-0.0234375,-0.0234375,0.0546875,0.015625,0.046875,0.03125,0.0859375,0.078125,0.078125,0.015625,-0.0234375,0.0390625,-0.03125,-0.046875,-0.0546875,0.015625,0.0234375,0.0,-0.0234375,-0.0078125,-0.015625,0.0078125,0.03125,-0.0,0.015625,-0.0390625,-0.015625,-0.0,-0.0078125,-0.0234375,-0.015625,-0.0078125,-0.0,-0.03125,-0.0,-0.0078125,0.015625,0.0,0.0234375,0.0234375,0.0859375,0.0,0.0859375,0.0,0.03125,-0.0390625,-0.0625,-0.078125,-0.046875,0.0,0.03125,-0.0078125,-0.078125,0.0234375,-0.0078125,0.03125,0.0703125,-0.0078125,-0.0390625,-0.0,0.015625,0.015625,-0.0078125,0.0078125,0.0234375,0.015625,-0.0078125,0.0,-0.0078125,-0.03125,-0.015625,-0.0234375,-0.0078125,0.015625,-0.0234375,0.0234375,-0.0390625,-0.0078125,-0.0625,0.015625,-0.0234375,0.0703125,-0.046875,-0.0234375,0.046875,-0.0078125,0.0625,0.015625,0.015625,-0.03125,-0.015625,0.0,0.015625,0.046875,-0.0234375,0.0234375,0.03125,0.046875,0.0390625,0.078125,-0.078125,0.0859375,0.0,0.0390625,0.015625,0.046875,-0.0546875,0.0078125,-0.0078125,-0.1171875,0.0234375,0.0234375,-0.03125,0.03125,0.0625,-0.0234375,0.078125,-0.0078125,-0.0078125,0.0234375,0.0078125,-0.0234375,0.03125,0.015625,-0.015625,-0.0390625,-0.0859375,0.1015625,-0.0546875,0.0625,-0.03125,0.046875,0.015625,0.0078125,-0.015625,-0.046875,-0.0859375,-0.0859375,-0.0546875,-0.0625,-0.015625,0.0234375,-0.0,0.0234375,0.0234375,0.015625,-0.0703125,-0.0390625,-0.09375,-0.0078125,0.0078125,-0.0078125,0.0,-0.0078125,-0.015625,0.0234375,-0.0390625,-0.03125,-0.1015625,0.046875,-0.0859375,0.03125,-0.0078125,-0.0390625,-0.0234375,-0.0390625,-0.015625,-0.0625,-0.015625,-0.015625,0.0078125,0.0,-0.0546875,0.0703125,0.0,0.0078125,0.1328125,0.0234375,0.0234375,0.046875,-0.0390625,0.0078125,0.0390625,-0.015625,-0.0703125,-0.03125,0.0234375,0.046875,0.03125,-0.015625,-0.0,-0.03125,-0.015625,-0.0625,0.0390625,0.078125,0.0078125,-0.0078125,-0.0703125,-0.0546875,-0.046875,-0.046875,-0.03125,-0.0625,0.0078125,-0.0390625,-0.03125,0.03125,-0.0234375,-0.0234375,0.140625,-0.046875,-0.0078125,0.0,-0.0078125,0.0,-0.0078125,0.0,-0.0078125,0.015625,0.0078125,0.0,-0.0078125,0.0078125,0.0546875,0.0390625,-0.0703125,0.0703125,0.0,-0.0390625,-0.046875,0.0546875,-0.0625,0.0234375,0.0703125,-0.0078125,0.0625,-0.0546875,-0.03125,-0.0546875,-0.015625,-0.0078125,0.0078125,-0.0625,-0.015625,-0.078125,0.0390625,0.109375,0.046875,-0.0078125,-0.0078125,-0.0078125,-0.0078125,0.0078125,0.0,0.0,0.0078125,-0.0078125,-0.0,0.0546875,0.046875,0.0859375,-0.015625,-0.046875,-0.0546875,0.03125,-0.015625,0.03125,0.0078125,-0.078125,-0.046875,-0.03125,-0.09375,0.0390625,0.015625,0.0390625,-0.0078125,-0.0546875,0.03125,0.0,0.015625,-0.0234375,-0.0078125,0.03125,0.0234375,-0.0234375,0.046875,-0.0234375,0.03125,0.0078125,0.0078125,0.03125,-0.0,0.03125,0.0078125,-0.046875,0.03125,-0.0625,-0.0234375,0.015625,-0.015625,-0.0078125,-0.03125,0.015625,0.0625,-0.015625,-0.0546875,-0.0,-0.0234375,-0.0390625,0.046875,0.0078125,-0.03125,0.046875,-0.015625,-0.03125,-0.03125,0.03125,-0.0078125,-0.0390625,-0.0,0.0078125,0.0390625,0.03125,0.0078125,-0.03125,-0.0234375,-0.0703125,0.015625,-0.0,0.03125,-0.015625,0.0078125,0.03125,0.03125,-0.0078125,0.0234375,-0.0546875,-0.03125,-0.0,-0.1171875,-0.0078125,-0.015625,-0.0,0.0546875,0.03125,0.0625,-0.0390625,0.0,0.0,-0.015625,-0.0,0.0078125,0.0078125,0.015625,0.0,0.0,0.0234375,0.0625,-0.0546875,0.0078125,-0.015625,0.0234375,-0.03125,-0.0625,0.0234375,-0.046875,0.0078125,-0.0625,-0.03125,0.015625,0.078125,0.0078125,0.0,0.015625,-0.0078125,-0.0546875,-0.0546875,-0.0234375,0.046875,-0.0,-0.0625,0.0390625,-0.0234375,-0.0703125,0.015625,0.0625,-0.0625,-0.03125,-0.0625,0.015625,0.0234375,0.109375,0.015625,0.0625,-0.03125,0.0,-0.03125,0.0390625,0.015625,0.015625,0.03125,0.015625,-0.0546875,0.09375,0.015625,0.0,0.015625,0.0078125,0.0,-0.015625,-0.0234375,-0.0390625,0.0,0.03125,-0.03125,0.125,0.015625,0.015625,-0.0859375,0.046875,0.0234375,0.03125,0.0078125,-0.03125,0.0390625,-0.0390625,-0.0234375,0.03125,0.0546875,0.0078125,0.015625,-0.046875,0.0703125,-0.0625,-0.0078125,-0.0078125,-0.0078125,-0.0078125,0.046875,0.046875,-0.0,-0.109375,-0.015625,0.0078125,0.015625,-0.046875,-0.1015625,0.125,-0.015625,-0.015625,-0.078125,0.0234375,0.0,0.0234375,0.03125,-0.046875,0.0390625,0.046875,0.0078125,0.03125,-0.0,-0.0546875,-0.03125,-0.03125,0.046875,0.0234375,-0.015625,0.046875,-0.03125,0.0546875,-0.0703125,-0.015625,-0.03125,-0.0078125,-0.078125,0.0546875,-0.0859375,-0.0078125,-0.0546875,0.0546875,0.0625,-0.0078125,-0.015625,-0.0078125,-0.0390625,-0.0390625,0.0546875,-0.0234375,-0.015625,0.0703125,0.0078125,0.015625,0.0703125,0.0,-0.0625,-0.0625,0.0078125,-0.0078125,-0.03125,-0.03125,0.0078125,0.0078125,-0.015625,0.0078125,0.015625,0.0,-0.0078125,-0.0,0.0078125,-0.0078125,-0.0234375,-0.046875,-0.0390625,0.0234375,-0.0390625,0.015625,0.0390625,-0.0390625,0.03125,0.0,-0.046875,-0.03125,-0.0625,-0.0625,0.015625,0.0234375,0.0078125,-0.0859375,0.0546875,-0.0234375,0.078125,0.0859375,-0.0625,0.0234375,-0.1015625,-0.0390625,0.0,0.0,-0.0078125,0.0,-0.0,-0.0078125,0.0078125,-0.015625,0.0,-0.0,-0.078125,-0.078125,0.109375,-0.015625,-0.0625,0.1015625,0.015625,0.0390625,-0.0234375,-0.078125,-0.0703125,0.015625,0.0078125,0.015625,0.046875,0.0,0.0234375,-0.09375,-0.0,-0.0234375,0.0,0.0546875,-0.0625,-0.0546875,-0.015625,-0.046875,0.046875,0.0,0.0,-0.046875,-0.0078125,-0.015625,-0.0234375,0.0390625,-0.046875,0.03125,-0.0078125,-0.03125,-0.03125,0.046875,-0.0,0.0078125,-0.015625,-0.046875,0.0546875,0.015625,-0.0390625,0.0078125,-0.03125,0.0234375,-0.0234375,-0.015625,0.046875,-0.0078125,-0.015625,0.0234375,0.0703125,0.03125,-0.03125,0.015625,0.015625,0.015625,0.0,0.03125,-0.0078125,0.0859375,0.0390625,0.015625,-0.0390625,-0.0078125,-0.0234375,0.015625,-0.046875,-0.0078125,-0.0859375,-0.0625,0.0234375,-0.0625,0.0234375,-0.0078125,-0.0078125,-0.046875,-0.0390625,0.0,0.0703125,-0.0625,0.0390625,-0.046875,-0.0234375,-0.0234375,-0.0234375,0.0078125,0.0234375,-0.0078125,-0.0,0.0078125,-0.0078125,-0.0078125,0.0234375,0.0546875,-0.0234375,-0.0390625,-0.0546875,0.0078125,-0.0078125,0.0390625,0.0234375,-0.0390625,-0.0078125,-0.046875,0.0234375,-0.0390625,0.0625,0.015625,0.0234375,0.03125,-0.0234375,-0.078125,-0.078125,-0.0234375,0.0625,0.0078125,-0.078125,-0.0859375,-0.078125,0.0234375,0.0625,-0.015625,0.0078125,-0.015625,0.0546875,0.0390625,-0.046875,0.015625,-0.0390625,-0.046875,-0.03125,0.0703125,-0.0234375,0.0546875,-0.0703125,-0.0546875,-0.0390625,-0.015625,0.0390625,-0.0078125,0.0078125,-0.046875,-0.046875,0.0,-0.0078125,0.015625,-0.0390625,0.015625,0.0234375,-0.015625,-0.1171875,0.0,0.0234375,-0.0625,0.03125,-0.03125,0.03125,-0.0234375,-0.0625,-0.0546875,0.0078125,0.015625,-0.0078125,-0.03125,0.0546875,0.0546875,0.09375,-0.0234375,-0.0546875,-0.046875,-0.046875,-0.0546875,-0.0625,-0.0546875,-0.0234375,-0.03125,0.078125,0.125,0.0078125,-0.0,-0.0,0.0390625,0.046875,0.015625,-0.0078125,0.1015625,0.0,-0.1015625,-0.0390625,-0.0,-0.0546875,0.0078125,0.0078125,-0.03125,-0.015625,-0.0546875,0.0390625,0.03125,-0.078125,-0.0390625,0.109375,0.0,0.015625,0.0546875,-0.0625,0.015625,0.0703125,-0.015625,-0.046875,0.015625,0.03125,-0.0078125,-0.0234375,0.015625,0.015625,0.015625,0.015625,-0.03125,0.015625,-0.0234375,0.015625,-0.0078125,-0.140625,0.03125,-0.0234375,-0.046875,0.0234375,-0.03125,-0.03125,-0.09375,0.015625,-0.0390625,-0.015625,-0.0625,0.0546875,0.0625,0.0,-0.0078125,-0.015625,0.0234375,0.0078125,-0.0078125,-0.015625,0.0078125,-0.0,0.0234375,0.015625,0.046875,0.0078125,-0.1171875,-0.078125,-0.015625,0.0546875,0.046875,0.015625,0.0390625,0.03125,0.0078125,-0.046875,-0.0234375,-0.0234375,-0.015625,0.0,0.0703125,0.0390625,-0.0703125,-0.046875,-0.0390625,0.09375,0.015625,-0.03125,-0.0390625,-0.0078125,-0.0078125,0.0078125,0.015625,-0.0,-0.0078125,0.0078125,0.0078125,-0.0,-0.0234375,-0.0859375,0.0234375,-0.03125,0.0234375,-0.03125,0.015625,-0.0,0.0703125,-0.0234375,0.1171875,0.015625,-0.0078125,-0.0625,-0.0234375,0.1015625,0.078125,0.1484375,0.03125,-0.0703125,0.0859375,-0.0,-0.1015625,-0.0546875,-0.0703125,0.1015625,0.0390625,0.0078125,0.0390625,-0.0,0.0234375,-0.046875,-0.015625,-0.0703125,0.0078125,-0.0,-0.0703125,-0.0234375,0.078125,-0.0234375,0.03125,0.0546875,-0.03125,0.0078125,0.0234375,0.0,-0.015625,0.0703125,0.03125,-0.0234375,0.09375,0.0,-0.015625,0.0078125,0.0390625,-0.0390625,0.078125,-0.0234375,-0.0546875,0.0234375,-0.0078125,0.0390625,0.03125,-0.0234375,-0.0546875,0.0,-0.0234375,-0.015625,0.015625,0.0078125,-0.046875,-0.046875,-0.0390625,0.0703125,-0.0078125,0.03125,-0.0078125,0.0078125,-0.0234375,-0.0546875,-0.0625,-0.0390625,0.0546875,-0.015625,-0.0234375,0.015625,-0.109375,0.0234375,-0.0390625,-0.0390625,-0.0,-0.0234375,-0.015625,-0.015625,0.0,-0.0,0.0078125,-0.0234375,-0.0078125,-0.0234375,0.0390625,0.1015625,-0.0234375,-0.015625,0.078125,-0.0390625,-0.078125,0.015625,-0.0546875,-0.015625,-0.03125,-0.0390625,-0.0234375,0.0390625,0.0234375,0.0234375,-0.0,-0.0078125,0.0390625,0.0078125,-0.046875,-0.078125,0.0546875,-0.0390625,-0.03125,0.0859375,-0.0078125,-0.015625,-0.0546875,-0.078125,-0.0703125,-0.046875,-0.0390625,-0.1015625,0.015625,0.0078125,-0.0234375,0.0546875,-0.0390625,0.0078125,0.0234375,-0.0546875,0.0234375,-0.0078125,-0.0078125,-0.0390625,0.0078125,0.0546875,-0.0625,0.0390625,0.1015625,0.0546875,0.0390625,-0.0859375,0.0625,-0.015625,0.0078125,-0.0703125,-0.0859375,0.1015625,-0.1171875,-0.0625,0.0234375,-0.0078125,-0.0390625,0.0234375,0.0390625,0.0,0.015625,-0.0390625,-0.03125,0.015625,-0.0078125,0.0,0.0234375,0.0625,0.0859375,0.109375,0.015625,0.0234375,0.03125,-0.0078125,0.0546875,-0.0625,0.0078125,0.0,-0.03125,-0.0234375,0.0390625,0.0859375,0.0390625,0.0703125,-0.078125,-0.046875,-0.09375,-0.0546875,0.03125,-0.0234375,0.0,0.0234375,0.0546875,-0.078125,-0.0859375,-0.09375,-0.1015625,0.03125,-0.0078125,0.0625,-0.046875,0.109375,-0.0,-0.09375,0.0625,0.0703125,0.046875,-0.03125,0.078125,0.015625,-0.0234375,-0.0078125,-0.0234375,-0.0390625,0.09375,0.015625,0.03125,0.0390625,0.0546875,-0.015625,-0.015625,0.0078125,-0.0390625,0.046875,-0.0234375,0.03125,0.078125,0.0078125,-0.0390625,-0.046875,0.0078125,0.0,0.046875,0.015625,-0.015625,-0.0078125,-0.0078125,0.0078125,-0.0,-0.0078125,-0.015625,-0.0,-0.0078125,-0.015625,-0.0625,0.03125,0.015625,-0.1015625,-0.0,0.0078125,0.03125,0.0546875,-0.0078125,-0.015625,-0.125,0.0078125,-0.03125,0.0546875,-0.0234375,-0.015625,0.0,-0.015625,0.078125,0.015625,-0.0078125,0.0390625,0.0390625,-0.0234375,-0.15625,-0.0625,-0.0078125,0.0078125,-0.0,-0.0,-0.0,-0.0078125,-0.0078125,0.0,-0.0078125,-0.0078125,0.0703125,-0.0078125,-0.0234375,0.015625,-0.046875,-0.015625,-0.0390625,0.0859375,-0.0390625,-0.0390625,-0.078125,-0.0,-0.015625,0.0078125,-0.03125,0.0625,-0.0078125,-0.0078125,-0.0234375,-0.0703125,-0.0078125,-0.0234375,0.0625,-0.015625,0.0234375,-0.078125,-0.015625,-0.0234375,-0.0078125,0.0078125,-0.0390625,-0.015625,0.0078125,0.0546875,-0.015625,0.0234375,-0.0,0.015625,0.0078125,0.078125,-0.0546875,-0.015625,0.0234375,0.0078125,-0.0390625,-0.0078125,-0.015625,-0.015625,-0.03125,-0.03125,-0.0078125,0.0078125,-0.03125,-0.015625,0.0390625,0.0078125,-0.0,-0.0,0.015625,-0.0078125,0.0078125,0.015625,0.0,-0.0078125,0.0078125,-0.0078125,-0.0625,0.0234375,-0.0,-0.046875,0.0078125,-0.015625,0.015625,-0.0,-0.03125,-0.0078125,0.0078125,-0.0078125,0.0078125,-0.0234375,-0.0234375,0.1015625,-0.015625,-0.0546875,-0.0234375,-0.0703125,-0.046875,-0.0390625,-0.0390625,-0.015625,-0.015625,-0.0078125,-0.0078125,-0.015625,0.0078125,-0.015625,0.0078125,-0.015625,-0.0,0.0078125,-0.015625,0.015625,-0.015625,-0.0234375,-0.0078125,0.0,0.0234375,0.0,-0.0078125,0.0234375,-0.0,-0.0078125,-0.0234375,-0.03125,0.0,0.015625,-0.0234375,-0.03125,0.0,0.015625,-0.0625,-0.0546875,-0.0234375,0.0078125,-0.015625,-0.0078125,0.0703125,0.015625,-0.0625,0.0234375,-0.0546875,-0.0546875,-0.015625,-0.0234375,-0.0078125,0.03125,-0.0234375,-0.0078125,0.0234375,-0.046875,-0.0078125,0.0859375,0.015625,0.0078125,-0.015625,0.0625,0.0078125,-0.046875,-0.015625,-0.0078125,-0.015625,0.0234375,-0.0078125,-0.0078125,0.0234375,-0.015625,-0.1171875,0.078125,-0.0234375,-0.109375,0.0078125,0.0,0.0390625,0.015625,-0.015625,0.015625,-0.0078125,0.0078125,0.015625,0.0390625,0.015625,-0.03125,0.0234375,-0.0078125,0.03125,-0.0078125,-0.0234375,-0.0625,0.0,-0.0,0.03125,0.015625,-0.015625,0.0390625,0.03125,-0.0390625,-0.03125,-0.0078125,0.0078125,0.015625,-0.0078125,-0.0546875,0.0625,0.03125,0.0078125,-0.0234375,-0.0625,-0.0234375,0.125,0.1015625,-0.0078125,0.046875,-0.0234375,-0.015625,0.015625,0.0,-0.0078125,-0.0234375,-0.03125,-0.015625,-0.015625,-0.015625,-0.015625,-0.03125,0.0234375,-0.03125,0.0,0.03125,-0.0078125,-0.0859375,-0.015625,-0.015625,0.0078125,-0.015625,-0.0078125,-0.0078125,0.0234375,-0.0234375,-0.015625,-0.0859375,-0.0546875,-0.0234375,0.0078125,-0.0078125,0.0703125,0.09375,0.078125,-0.0390625,-0.0390625,0.015625,-0.0078125,-0.03125,-0.0078125,0.0078125,-0.0078125,0.0,-0.0078125,-0.015625,0.0078125,-0.0078125,0.015625,0.015625,0.015625,0.078125,-0.015625,-0.015625,-0.0703125,-0.09375,-0.0,0.0546875,0.109375,-0.0234375,-0.015625,0.0625,-0.0234375,0.03125,-0.0390625,0.0234375,-0.0078125,-0.0234375,0.0078125,0.0234375,-0.0078125,0.078125,-0.0078125,0.078125,-0.015625,-0.03125,-0.015625,-0.0,0.0,0.0078125,0.0,-0.0078125,0.0078125,-0.0078125,0.0078125,0.0078125,0.015625,-0.015625,-0.0078125,-0.0078125,-0.0625,-0.09375,-0.0390625,0.0234375,-0.0078125,0.0234375,0.0078125,0.0625,-0.0390625,-0.0234375,0.03125,-0.0390625,-0.015625,0.03125,-0.0234375,0.046875,-0.03125,-0.015625,0.03125,-0.0078125,-0.015625,-0.046875,-0.0703125,0.03125,0.0078125,-0.0078125,-0.0390625,0.015625,-0.0234375,-0.0234375,-0.0234375,0.0234375,0.0234375,-0.046875,-0.0234375,-0.0546875,0.0078125,-0.0390625,-0.0234375,0.015625,-0.0703125,0.0078125,0.0078125,0.0546875,0.0,-0.015625,0.0,-0.015625,0.03125,0.0234375,0.0,0.03125,-0.0078125,-0.0078125,0.0234375,0.015625,-0.0234375,-0.0234375,0.0234375,-0.015625,-0.0234375,-0.0234375,-0.015625,0.0078125,-0.0078125,-0.015625,-0.0625,0.0234375,0.1640625,-0.046875,0.125,-0.046875,-0.0703125,-0.078125,-0.0078125,-0.0625,0.015625,0.0078125,-0.046875,0.03125,-0.015625,-0.015625,0.0390625,-0.03125,0.046875,-0.0625,0.0234375,0.0078125,0.0078125,-0.0078125,-0.0,0.0,-0.0,0.0,-0.0234375,-0.0390625,-0.015625,-0.0234375,-0.015625,0.0234375,-0.0390625,-0.015625,0.0390625,0.0078125,0.09375,-0.015625,0.0078125,0.015625,0.0390625,-0.0234375,-0.0390625,-0.046875,0.03125,-0.0078125,0.0078125,-0.0625,-0.0234375,-0.1015625,-0.0625,-0.046875,0.0234375,0.125,0.03125,-0.03125,-0.0625,0.0390625,-0.0078125,0.09375,-0.0234375,-0.046875,0.0,0.046875,0.015625,-0.0078125,-0.03125,0.03125,-0.03125,-0.0390625,0.046875,0.0,0.078125,0.03125,0.0625,-0.015625,-0.0703125,-0.0234375,-0.0078125,0.0390625,-0.0234375,-0.0546875,-0.0546875,-0.0234375,-0.0078125,0.0078125,-0.03125,-0.0390625,0.0,0.15625,-0.0390625,0.015625,-0.0625,-0.0390625,-0.0078125,-0.015625,-0.03125,0.03125,0.1015625,0.0390625,0.03125,-0.0234375,0.0078125,-0.0546875,-0.0,-0.03125,-0.0078125,-0.0390625,0.0,0.046875,0.03125,-0.0234375,0.0078125,-0.0,-0.0390625,-0.0234375,-0.0390625,0.0078125,-0.1875,0.0078125,-0.0234375,0.0234375,0.0390625,-0.046875,-0.0078125,-0.015625,0.0546875,-0.0546875,0.03125,-0.046875,-0.0234375,-0.015625,0.0234375,-0.0234375,-0.0078125,0.0546875,-0.03125,0.03125,-0.03125,-0.0703125,-0.0859375,-0.015625,0.0078125,-0.046875,0.03125,-0.1015625,-0.0390625,0.0078125,-0.015625,0.0390625,-0.0078125,0.0703125,0.0546875,-0.046875,0.0078125,0.0390625,0.015625,0.0390625,-0.0,-0.0390625,-0.078125,-0.03125,-0.015625,-0.015625,0.03125,-0.046875,-0.0390625,0.0078125,-0.0703125,-0.0390625,-0.0546875,0.0078125,0.015625,0.0078125,-0.015625,0.0234375,-0.0078125,-0.0078125,0.0078125,-0.0078125,-0.0234375,-0.0234375,-0.0234375,-0.0,-0.046875,0.0078125,0.03125,-0.0234375,-0.03125,-0.0078125,0.0078125,0.0,-0.0234375,-0.046875,-0.0390625,0.046875,0.0234375,-0.0078125,-0.0,-0.015625,-0.0078125,-0.046875,0.0078125,-0.0546875,-0.0,0.171875,0.03125,-0.0078125,0.0,-0.0078125,0.0078125,0.0078125,0.0078125,0.015625,0.0078125,0.0078125,-0.0,-0.03125,-0.0234375,0.046875,-0.03125,-0.1015625,0.0703125,0.046875,-0.0390625,0.0,-0.0546875,0.0,-0.046875,-0.0078125,-0.0625,0.03125,0.046875,-0.0078125,-0.0234375,-0.015625,-0.0078125,-0.0234375,-0.1328125,-0.078125,-0.03125,0.09375,0.0234375,-0.015625,-0.0390625,-0.03125,-0.0390625,0.03125,-0.0234375,-0.0,-0.0625,0.0390625,-0.0234375,-0.0078125,0.015625,-0.0234375,-0.015625,-0.046875,0.0234375,0.0390625,-0.0390625,0.0,-0.0078125,0.0078125,-0.0625,0.09375,0.03125,-0.0078125,0.0078125,-0.015625,0.0390625,0.0078125,-0.015625,-0.0,-0.0703125,0.0390625,0.015625,0.03125,-0.0234375,0.0,-0.0078125,-0.0078125,0.0078125,-0.046875,-0.015625,-0.046875,-0.0234375,-0.0234375,-0.0234375,-0.015625,-0.015625,-0.0859375,0.046875,-0.0859375,-0.0546875,0.03125,-0.0,-0.0390625,-0.015625,-0.0078125,-0.0390625,0.0390625,0.0390625,0.0078125,0.0078125,0.03125,0.0,-0.0,-0.0078125,-0.0,-0.0078125,0.0,-0.0234375,0.015625,-0.0078125,-0.015625,0.0078125,-0.015625,-0.015625,-0.0,-0.0,-0.015625,-0.0390625,-0.0078125,-0.015625,-0.0234375,-0.015625,0.03125,0.0390625,0.140625,-0.046875,0.0,0.0625,-0.015625,0.0,0.0078125,-0.0234375,0.0390625,0.03125,0.0234375,0.0625,-0.0625,0.0,-0.0390625,0.0078125,-0.015625,0.0703125,-0.015625,-0.0390625,-0.0390625,-0.0234375,-0.0,-0.03125,-0.015625,-0.0625,0.0,-0.015625,-0.0,-0.09375,0.015625,0.0078125,-0.0078125,0.0,-0.0546875,-0.0234375,-0.015625,-0.078125,0.015625,-0.0390625,-0.015625,-0.015625,-0.015625,-0.0234375,-0.09375,0.03125,-0.0234375,-0.0703125,0.015625,-0.0390625,-0.0234375,-0.015625,-0.0078125,0.0546875,-0.0859375,-0.015625,0.0390625,0.046875,0.0234375,-0.0078125,0.015625,-0.0390625,-0.0390625,-0.0234375,-0.0859375,0.1328125,-0.0078125,0.03125,0.0390625,0.0,0.0234375,-0.1328125,-0.015625,-0.0390625,-0.015625,-0.0546875,-0.0,-0.0078125,-0.03125,-0.0234375,-0.03125,-0.03125,0.1015625,-0.046875,0.0625,-0.0078125,0.0078125,-0.0078125,0.046875,0.03125,0.0078125,0.03125,-0.03125,-0.078125,0.03125,0.03125,-0.0234375,0.0078125,-0.09375,0.0703125,0.0234375,-0.0625,-0.0546875,0.0390625,-0.0,0.015625,0.0546875,-0.078125,-0.0546875,-0.015625,0.015625,-0.0078125,-0.0,-0.015625,-0.015625,-0.0546875,0.0390625,0.1171875,-0.0078125,-0.0625,-0.046875,-0.03125,0.03125,0.125,-0.015625,-0.0234375,-0.0,0.0078125,-0.0234375,-0.0078125,-0.0078125,-0.0078125,0.015625,-0.0078125,-0.015625,-0.015625,-0.0,-0.0078125,-0.0078125,0.0,-0.09375,-0.09375,-0.0,-0.0078125,-0.0078125,-0.0,0.015625,0.0,-0.03125,-0.0703125,-0.03125,-0.015625,0.046875,-0.0078125,-0.015625,0.0234375,0.0,-0.0078125,-0.0390625,-0.015625,-0.0078125,-0.0390625,-0.109375,0.0078125,-0.0546875,0.03125,-0.0078125,0.0078125,0.015625,-0.015625,0.0,-0.015625,-0.0078125,0.0,0.0,-0.015625,-0.0234375,0.0234375,-0.0078125,-0.0,-0.03125,-0.015625,-0.015625,-0.03125,-0.0078125,0.0625,0.078125,-0.03125,-0.03125,-0.0234375,0.0,0.0078125,0.0078125,0.015625,0.046875,0.0390625,-0.03125,-0.09375,0.03125,0.0078125,-0.03125,0.0234375,-0.015625,-0.078125,0.0078125,-0.0234375,0.0234375,0.0703125,0.015625,0.0234375,0.0078125,-0.0234375,-0.0234375,0.0859375,0.0,-0.0078125,-0.0078125,0.0,0.0,-0.0703125,0.0,0.0078125,0.0,-0.0078125,0.0,0.03125,-0.015625,-0.0078125,-0.0078125,0.0078125,0.0078125,0.0,0.0078125,-0.0,0.0234375,-0.0078125,0.015625,-0.0078125,-0.015625,-0.015625,-0.0078125,-0.0,0.015625,0.0078125,-0.03125,0.0390625,0.046875,0.0,-0.0,0.0078125,-0.0,0.046875,-0.0625,0.03125,0.0390625,-0.0078125,0.03125,-0.046875,-0.0390625,0.0078125,-0.046875,0.046875,0.0234375,-0.03125,-0.046875,-0.0,-0.0078125,-0.015625,-0.0,0.0078125,-0.015625,0.0078125,-0.0078125,0.015625,-0.0234375,-0.015625,0.015625,-0.03125,-0.0,0.0,-0.03125,-0.0390625,-0.0234375,-0.015625,-0.03125,-0.0625,-0.015625,0.0625,-0.0234375,0.015625,0.109375,-0.03125,-0.0,0.03125,-0.03125,-0.0234375,-0.046875,-0.0546875,0.03125,0.0625,0.0546875,-0.0078125,0.0390625,-0.125,-0.0078125,0.03125,-0.125,0.0,0.0234375,0.0859375,-0.0234375,0.03125,0.0078125,-0.015625,-0.0234375,-0.0234375,0.0078125,-0.046875,0.0078125,-0.0234375,0.046875,-0.0390625,0.0234375,-0.0234375,-0.078125,0.0234375,-0.015625,0.0234375,-0.015625,0.03125,-0.0546875,-0.0078125,0.0390625,0.1640625,-0.0234375,0.09375,-0.0625,-0.0078125,-0.015625,0.0390625,-0.015625,-0.03125,-0.0234375,-0.0078125,-0.046875,-0.0546875,-0.0078125,-0.046875,0.046875,-0.0234375,0.0234375,-0.0390625,-0.03125,0.03125,-0.0234375,-0.0,0.046875,0.0234375,-0.015625,0.015625,-0.0625,0.0078125,-0.0703125,0.0859375,0.015625,0.0390625,-0.0625,0.0,-0.0703125,0.0390625,-0.0390625,-0.03125,-0.0390625,-0.0390625,-0.015625,-0.0078125,-0.0390625,-0.0390625,-0.109375,-0.0078125,0.015625,0.09375,-0.0234375,-0.0625,-0.0078125,-0.03125,0.0703125,-0.0,-0.0078125,-0.0546875,-0.03125,-0.03125,0.0,0.0390625,-0.015625,-0.046875,-0.0546875,0.0078125,0.0078125,-0.0546875,-0.0078125,0.109375,0.1484375,-0.015625,-0.0390625,0.03125,0.0,-0.0390625,-0.0390625,0.015625,-0.0546875,0.0078125,0.078125,0.0078125,-0.0390625,-0.046875,-0.078125,-0.015625,0.0078125,0.0,0.0078125,0.0078125,-0.0078125,-0.0,0.0078125,-0.015625,0.0,-0.046875,0.0390625,0.0078125,-0.0390625,-0.0703125,-0.0078125,0.0390625,-0.0703125,-0.0234375,0.0234375,-0.0234375,0.015625,0.0390625,-0.0390625,0.015625,0.0625,-0.0546875,0.0078125,0.0,-0.0234375,-0.0390625,0.015625,-0.0,-0.0078125,-0.03125,0.0546875,0.015625,0.0,-0.0078125,0.0078125,0.0078125,0.0,0.0,0.0078125,-0.0078125,-0.0078125,0.015625,-0.0390625,-0.0234375,-0.0078125,0.03125,-0.0390625,-0.0234375,0.015625,-0.0,-0.0859375,0.03125,0.03125,0.0859375,-0.0625,-0.015625,0.0078125,-0.078125,-0.015625,0.0625,-0.0234375,0.0234375,0.015625,-0.0078125,0.015625,-0.0625,0.0234375,-0.0234375,-0.0234375,0.0390625,0.03125,0.015625,-0.0390625,-0.0078125,0.046875,0.0078125,0.0078125,0.0,-0.015625,-0.0078125,-0.03125,-0.0234375,-0.0078125,0.015625,-0.0703125,0.015625,0.0078125,0.015625,0.015625,-0.0625,-0.03125,-0.0234375,0.03125,-0.03125,0.0234375,-0.0,0.0078125,0.0234375,-0.0,0.0,0.0,0.0078125,-0.0234375,-0.015625,0.0078125,-0.015625,-0.015625,-0.0234375,0.0234375,0.0,0.0546875,-0.03125,-0.015625,0.078125,-0.03125,-0.0078125,-0.078125,-0.0859375,0.0234375,0.0546875,-0.109375,-0.0078125,-0.03125,0.0078125,0.015625,-0.0,0.09375,-0.03125,-0.109375,0.0078125,0.015625,-0.015625,0.0078125,0.015625,-0.015625,-0.0078125,-0.0078125,0.0,0.0,-0.0,-0.046875,-0.03125,0.0078125,-0.015625,-0.0078125,-0.0078125,-0.015625,-0.015625,-0.0234375,0.015625,-0.0,0.0078125,-0.015625,-0.0390625,-0.046875,0.1171875,-0.0703125,-0.015625,0.0078125,-0.03125,-0.03125,0.171875,-0.0546875,0.0078125,0.1640625,-0.0625,-0.0078125,0.0390625,0.0078125,0.0390625,-0.1015625,-0.015625,-0.03125,0.046875,0.03125,-0.0234375,0.0078125,-0.015625,0.0859375,-0.046875,-0.0078125,0.0,0.0078125,0.0390625,0.015625,0.0390625,0.0390625,-0.0390625,-0.0625,0.046875,-0.0390625,-0.0234375,-0.0546875,-0.0078125,-0.046875,-0.0390625,0.0078125,0.0390625,0.0234375,0.0,0.1015625,-0.09375,-0.0234375,0.0078125,0.0078125,-0.0234375,0.0625,0.0078125,-0.0234375,-0.0078125,0.015625,-0.0078125,-0.015625,0.09375,-0.0078125,-0.1171875,-0.0078125,-0.015625,-0.0390625,-0.0625,-0.046875,-0.0859375,0.03125,0.0234375,0.0078125,-0.078125,-0.015625,-0.046875,0.015625,0.015625,0.015625,0.015625,-0.0390625,-0.0546875,-0.046875,-0.0234375,0.125,-0.0078125,-0.0625,-0.03125,-0.03125,-0.0234375,-0.03125,-0.0625,0.0078125,0.1015625,-0.0,0.0078125,-0.0625,0.046875,0.0078125,-0.078125,-0.0,0.015625,0.0234375,-0.0078125,-0.0390625,0.0390625,0.0625,-0.015625,-0.0703125,-0.0078125,-0.015625,-0.0,-0.03125,0.0078125,-0.0078125,0.0,0.0078125,0.09375,0.0234375,-0.03125,-0.046875,-0.0625,-0.0078125,-0.0390625,0.03125,0.1328125,-0.0078125,-0.0234375,0.0234375,0.0,-0.015625,-0.015625,-0.0,0.0078125,0.0078125,-0.0078125,-0.0078125,0.015625,-0.0,0.0078125,0.0,0.0234375,0.0390625,-0.0625,0.046875,0.0234375,-0.0078125,-0.015625,-0.015625,-0.0078125,-0.046875,0.046875,-0.015625,-0.046875,0.1015625,0.0234375,-0.0,-0.015625,-0.03125,0.03125,-0.0625,-0.0078125,0.0078125,-0.0234375,0.0625,-0.0078125,0.0390625,0.0,-0.0078125,0.0078125,0.0,-0.015625,0.0078125,-0.0,-0.015625,-0.0078125,-0.015625,-0.0078125,0.0703125,0.0,0.0078125,-0.03125,-0.03125,-0.0078125,0.0078125,0.0390625,-0.0390625,-0.0078125,-0.015625,-0.0625,-0.03125,0.078125,-0.0078125,0.015625,0.0,0.0078125,-0.0078125,0.015625,0.015625,0.015625,-0.03125,-0.0390625,-0.0546875,-0.046875,0.015625,-0.015625,0.0078125,0.0,-0.078125,0.0,-0.015625,-0.03125,-0.0390625,-0.03125,0.0,-0.0078125,-0.046875,0.0234375,0.0078125,-0.0078125,-0.0390625,0.03125,-0.0078125,0.015625,0.046875,-0.0078125,0.0,0.0390625,-0.0,0.0234375,-0.015625,-0.0234375,0.0078125,-0.0546875,-0.015625,-0.0078125,-0.0078125,0.0078125,-0.0078125,-0.0078125,0.0390625,-0.015625,-0.0390625,-0.046875,0.0625,0.0234375,-0.0,-0.0234375,0.03125,0.0078125,-0.078125,0.046875,-0.0078125,0.0078125,0.0234375,0.0,-0.0546875,-0.0078125,0.046875,0.03125,0.0,0.03125,0.0078125,-0.0703125,-0.03125,-0.015625,0.0234375,-0.0,0.0,-0.0078125,0.0078125,0.015625,0.015625,-0.0,0.0078125,0.0234375,-0.015625,-0.0078125,-0.015625,-0.0078125,-0.0390625,-0.03125,-0.0234375,0.0078125,-0.0078125,-0.03125,0.015625,0.0078125,-0.0234375,0.078125,-0.046875,-0.0,-0.0234375,0.0078125,0.0078125,-0.03125,0.0859375,0.0390625,-0.0078125,0.0234375,-0.03125,0.0078125,-0.046875,0.015625,-0.0546875,0.0703125,-0.0390625,-0.109375,-0.1015625,0.03125,0.03125,0.0078125,0.0,-0.0625,-0.0078125,0.0078125,0.015625,0.0,-0.0078125,0.0390625,-0.015625,-0.0234375,0.0234375,-0.0078125,0.0078125,-0.0078125,-0.0234375,-0.015625,-0.0,0.0,-0.0078125,0.0234375,0.015625,0.015625,-0.0703125,-0.015625,-0.046875,-0.015625,-0.0390625,-0.0625,0.0546875,-0.0078125,-0.0078125,-0.015625,0.0625,-0.0078125,0.0234375,-0.0234375,0.0,-0.0546875,-0.078125,0.0,0.0234375,0.0390625,0.0078125,-0.0,0.046875,-0.0,0.0078125,-0.03125,0.0234375,-0.03125,0.0,0.0078125,0.0234375,0.0234375,0.03125,0.0703125,-0.046875,-0.0078125,0.015625,-0.1015625,0.03125,-0.03125,0.0,0.0078125,-0.046875,-0.09375,-0.03125,0.015625,-0.0,0.0078125,-0.046875,0.078125,0.0625,-0.015625,-0.046875,-0.03125,0.015625,0.0,-0.015625,-0.1015625,0.03125,0.0546875,-0.1015625,-0.0078125,-0.0078125,-0.0625,-0.015625,0.0,-0.015625,-0.015625,-0.0078125,0.0546875,-0.0,-0.046875,-0.046875,-0.0078125,-0.03125,-0.046875,-0.015625,-0.0234375,0.0078125,0.0546875,-0.0390625,-0.0703125,0.0234375,0.0078125,0.0078125,0.0546875,0.0,-0.0078125,-0.0078125,-0.0078125,-0.0078125,-0.0078125,-0.0,0.0,0.0,-0.0234375,0.0546875,0.09375,0.03125,-0.0234375,-0.109375,-0.0078125,0.0078125,-0.0078125,-0.015625,0.0078125,0.0078125,-0.015625,0.0546875,-0.078125,0.0078125,-0.0546875,-0.0,0.046875,0.046875,-0.0234375,-0.03125,-0.0078125,-0.1328125,-0.078125,-0.03125,0.0078125,0.0078125,0.0078125,0.0234375,-0.0,0.0078125,0.0,0.0,-0.0078125,-0.015625,-0.015625,0.0078125,-0.0703125,0.078125,0.0703125,-0.0078125,-0.015625,-0.1015625,-0.03125,-0.0390625,-0.0390625,-0.046875,-0.046875,-0.0625,-0.0078125,-0.015625,0.03125,0.1171875,-0.0078125,0.03125,0.03125,0.015625,-0.03125,-0.078125,-0.0234375,0.046875,0.0390625,-0.015625,-0.03125,-0.015625,0.046875,-0.0703125,-0.125,0.03125,0.0390625,0.1015625,0.0234375,0.0078125,-0.0234375,-0.0,-0.0859375,-0.0234375,0.0078125,0.03125,-0.0625,-0.0,0.0234375,-0.046875,-0.0078125,0.0234375,0.0703125,-0.015625,0.0078125,0.03125,-0.015625,0.0078125,0.015625,0.0078125,0.0,0.09375,-0.015625,0.0,-0.0,0.0,-0.0078125,0.0703125,0.0234375,-0.0078125,-0.0546875,-0.046875,-0.03125,-0.046875,-0.015625,0.03125,-0.0703125,-0.03125,-0.015625,-0.0625,-0.0078125,0.0859375,0.0390625,0.0234375,-0.0,-0.0546875,0.0078125,0.0078125,-0.0,0.0078125,0.0,0.0625,-0.015625,-0.0078125,-0.0078125,-0.0078125,-0.0390625,-0.0078125,0.0078125,0.0078125,0.015625,-0.015625,0.03125,-0.0390625,0.0,-0.03125,0.0234375,0.0390625,-0.0546875,0.03125,0.0078125,-0.0546875,0.0234375,-0.015625,-0.046875,0.03125,-0.0078125,-0.0546875,0.0234375,-0.0078125,-0.015625,-0.0390625,-0.046875,0.03125,-0.078125,0.0,0.078125,0.0,0.0234375,-0.046875,0.125,0.0078125,-0.1171875,0.0,-0.0625,-0.046875,0.046875,-0.0234375,0.0546875,-0.1171875,-0.03125,-0.0234375,-0.0390625,-0.03125,0.046875,0.09375,0.015625,-0.046875,0.046875,-0.03125,-0.0,-0.0234375,0.015625,0.046875,-0.0234375,-0.0,0.0234375,0.0234375,-0.0078125,-0.0546875,-0.0234375,-0.0625,0.0234375,-0.0078125,0.0078125,0.0390625,-0.0703125,-0.03125,-0.015625,-0.0546875,0.0078125,0.0,0.125,0.0390625,-0.0546875,-0.0,0.0,-0.03125,0.03125,-0.015625,0.03125,0.0546875,-0.0234375,-0.015625,0.125,-0.0078125,-0.0234375,-0.0546875,-0.0234375,0.0625,0.0625,-0.03125,0.015625,0.0234375,0.015625,-0.0546875,0.140625,0.0234375,-0.078125,0.0234375,0.0625,-0.03125,0.1171875,0.0078125,-0.046875,0.0234375,-0.0703125,-0.0234375,-0.1015625,0.03125,0.0234375,0.03125,0.03125,-0.015625,-0.1171875,-0.015625,0.046875,-0.125,0.0703125,-0.0390625,0.109375,-0.0078125,-0.125,-0.109375,0.0078125,0.0234375,-0.0546875,0.015625,0.0390625,-0.0625,0.0234375,-0.03125,0.0078125,-0.015625,-0.0390625,-0.0625,-0.0390625,-0.0625,-0.015625,-0.015625,0.0859375,0.09375,0.0078125,-0.078125,-0.046875,0.0,-0.015625,-0.0078125,-0.0078125,-0.0078125,0.0,-0.015625,0.0,0.0078125,0.015625,0.0546875,-0.0078125,-0.0078125,-0.0859375,-0.03125,-0.0078125,0.0234375,-0.046875,0.015625,-0.0,-0.015625,0.015625,0.0625,-0.03125,-0.0390625,0.015625,-0.0078125,0.0078125,-0.0,0.0078125,0.0234375,0.0703125,-0.0546875,-0.0078125,-0.03125,-0.03125,-0.0078125,-0.015625,0.0078125,-0.0078125,-0.0,0.0078125,-0.0078125,0.0078125,-0.0,-0.015625,0.0234375,0.0,0.0,0.03125,-0.078125,-0.015625,-0.046875,-0.046875,0.0234375,0.0546875,-0.0625,-0.0078125,-0.0859375,-0.0703125,0.0390625,0.0390625,0.015625,-0.03125,0.0625,-0.015625,0.015625,0.015625,-0.046875,0.0234375,0.0078125,-0.046875,-0.015625,-0.03125,0.0234375,0.0,-0.0078125,-0.0390625,-0.0078125,-0.0078125,-0.0078125,-0.0390625,-0.0,0.015625,0.0,-0.046875,-0.0,0.0078125,-0.0546875,-0.0859375,-0.015625,-0.0234375,0.0,-0.015625,-0.015625,0.0390625,-0.015625,-0.0078125,0.0,0.015625,0.0234375,-0.0078125,-0.015625,-0.0078125,0.015625,-0.0078125,-0.0078125,0.046875,0.0234375,0.0390625,0.03125,-0.0078125,-0.0390625,-0.0078125,-0.0234375,-0.0390625,-0.09375,-0.0390625,-0.015625,-0.046875,0.015625,0.078125,-0.0703125,-0.0234375,-0.0,-0.0078125,0.0,0.0,-0.03125,-0.015625,-0.015625,0.0390625,-0.0234375,-0.0234375,0.1015625,-0.0,-0.0078125,-0.0,-0.0078125,0.0078125,-0.0,-0.0078125,-0.0,-0.015625,0.0390625,0.0,-0.0078125,-0.0078125,-0.046875,0.0234375,-0.0234375,0.015625,-0.0078125,0.015625,-0.0390625,-0.015625,-0.015625,-0.0234375,-0.0078125,0.0078125,-0.0546875,-0.0390625,-0.015625,-0.0078125,-0.0625,-0.03125,0.0625,0.0234375,-0.015625,-0.046875,-0.0859375,0.0078125,-0.078125,0.03125,-0.015625,-0.03125,0.1171875,-0.0390625,0.0,-0.0390625,0.0234375,-0.046875,-0.0390625,-0.0390625,0.0390625,-0.1015625,-0.0390625,-0.0,0.1171875,-0.03125,-0.0390625,0.03125,-0.0234375,-0.0234375,0.0546875,-0.0390625,-0.0078125,-0.046875,0.0078125,-0.015625,-0.0078125,-0.0234375,-0.015625,0.0546875,-0.015625,-0.015625,-0.046875,-0.0078125,-0.0546875,-0.0078125,0.015625,-0.0625,-0.0078125,-0.0078125,0.03125,-0.0,0.015625,-0.046875,0.046875,-0.046875,-0.109375,-0.0078125,-0.0234375,-0.0234375,0.0078125,0.0625,0.0625,-0.0234375,-0.0390625,0.0546875,0.015625,0.0078125,-0.046875,0.046875,0.0078125,-0.0078125,-0.1171875,-0.03125,-0.0078125,0.0703125,-0.0078125,-0.0234375,0.171875,0.0078125,-0.015625,0.0078125,-0.015625,-0.03125,0.015625,-0.0,-0.03125,-0.046875,0.015625,0.0078125,-0.046875,-0.046875,-0.0703125,-0.109375,0.0,0.125,-0.1484375,-0.0078125,0.03125,0.046875,-0.015625,-0.078125,0.125,-0.0390625,-0.03125,-0.109375,-0.0,-0.0546875,0.0390625,-0.0390625,0.0859375,-0.0234375,0.015625,-0.0078125,0.0,0.046875,-0.0234375,-0.0078125,0.0078125,-0.0234375,0.0078125,-0.015625,-0.0234375,0.046875,0.0078125,0.0078125,-0.0078125,-0.0078125,0.015625,-0.0078125,-0.0,0.0,0.0078125,0.015625,-0.03125,0.015625,-0.015625,-0.0,-0.015625,-0.046875,0.046875,0.0234375,0.0703125,-0.03125,-0.0234375,-0.0390625,-0.0390625,0.1171875,-0.0546875,-0.078125,0.0390625,-0.0703125,0.078125,-0.0078125,-0.0390625,-0.0078125,-0.0234375,-0.015625,0.0234375,-0.03125,-0.0078125,0.0078125,-0.015625,-0.0,0.0078125,-0.0078125,0.0078125,-0.0078125,0.0078125,0.1015625,0.0234375,0.0234375,0.0625,-0.0234375,-0.0390625,-0.046875,-0.015625,-0.0546875,0.0703125,0.0,-0.03125,0.03125,-0.015625,0.03125,-0.03125,0.0703125,-0.0078125,0.0078125,-0.046875,0.015625,-0.1015625,-0.09375,0.0390625,0.0546875,-0.0625,-0.0234375,0.015625,0.0234375,-0.0078125,-0.03125,-0.03125,0.0078125,0.0625,0.1015625,0.046875,0.046875,0.0703125,0.0546875,0.046875,-0.03125,-0.0390625,-0.015625,0.0390625,-0.03125,-0.0078125,-0.03125,0.03125,0.0390625,0.0703125,0.03125,-0.0234375,-0.0390625,-0.015625,-0.046875,-0.0546875,-0.03125,0.015625,0.046875,-0.0078125,-0.015625,0.015625,0.0078125,0.0078125,-0.015625,-0.0234375,0.0625,-0.015625,-0.0078125,-0.0390625,-0.046875,-0.0234375,0.0625,0.0859375,-0.0078125,-0.0703125,-0.046875,-0.0703125,-0.0,0.0390625,0.0625,0.015625,0.03125,0.0859375,-0.0078125,-0.0703125,-0.0625,0.0,-0.0,0.015625,0.0078125,0.0,0.0078125,0.015625,0.015625,0.0078125,0.0078125,-0.0078125,-0.0078125,0.0234375,-0.0078125,-0.0546875,0.0390625,-0.03125,0.046875,-0.0390625,0.0078125,0.03125,0.0078125,-0.0546875,-0.0390625,-0.0703125,-0.0625,-0.03125,0.0625,-0.046875,-0.0234375,-0.0078125,0.0546875,-0.0,-0.0859375,0.015625,-0.0234375,-0.0234375,0.03125,-0.0859375,0.03125,0.0859375,0.0390625,0.0078125,-0.0078125,-0.0703125,-0.0234375,0.015625,0.0078125,-0.046875,0.0078125,-0.09375,-0.0078125,0.0390625,-0.0703125,0.0078125,0.046875,0.0703125,-0.0234375,-0.015625,0.015625,0.0234375,-0.0625,-0.015625,-0.015625,-0.0390625,0.0078125,-0.0859375,0.0625,0.09375,-0.078125,-0.03125,-0.046875,-0.046875,0.0234375,-0.0703125,0.0078125,0.0234375,-0.03125,-0.015625,-0.0,-0.0234375,-0.0390625,-0.0078125,-0.03125,-0.0703125,-0.078125,0.0234375,-0.046875,-0.1015625,0.0,0.0,0.0078125,0.046875,-0.03125,-0.0625,-0.03125,-0.0,-0.015625,0.0859375,-0.0859375,-0.046875,-0.0234375,-0.046875,0.0078125,0.03125,-0.015625,-0.0703125,-0.046875,-0.03125,-0.015625,0.0234375,-0.0,0.078125,-0.0,-0.03125,0.1015625,-0.0,-0.0078125,0.0234375,-0.0546875,0.0546875,-0.0078125,0.015625,0.0859375,-0.0234375,-0.0234375,-0.0390625,-0.0078125,0.0,0.0390625,-0.03125,0.0390625,0.0078125,0.03125,-0.09375,-0.0234375,0.03125,-0.0,-0.078125,-0.0078125,0.046875,0.125,-0.0625,0.015625,0.015625,0.0078125,0.046875,0.0234375,-0.0078125,0.015625,-0.015625,-0.0,0.0625,-0.0703125,-0.0703125,0.0,-0.0078125,-0.0078125,0.0078125,0.015625,-0.015625,-0.015625,-0.015625,-0.0078125,-0.015625,-0.0,-0.0390625,-0.046875,-0.09375,-0.109375,0.015625,0.0546875,0.0078125,-0.015625,0.015625,-0.078125,-0.03125,-0.015625,-0.015625,-0.0234375,-0.046875,-0.0390625,-0.0234375,-0.03125,-0.015625,-0.015625,0.015625,-0.03125,-0.015625,0.125,-0.03125,-0.0234375,0.0078125,-0.0078125,0.0,0.0,0.0078125,-0.0078125,0.0078125,-0.0,0.0078125,-0.046875,-0.09375,-0.03125,-0.078125,0.03125,-0.0078125,-0.09375,0.125,-0.0,-0.109375,0.0390625,-0.0078125,0.0078125,-0.0,0.015625,-0.0859375,0.0,-0.0,0.03125,-0.0078125,-0.0078125,0.1015625,-0.0859375,-0.0390625,0.0859375,-0.078125,-0.0390625,0.046875,-0.0234375,0.015625,-0.0234375,0.0234375,0.0078125,0.0078125,0.015625,0.0,-0.0,0.0390625,-0.0390625,0.0234375,-0.015625,0.0078125,0.0,-0.0546875,-0.0078125,-0.0703125,-0.0234375,0.015625,-0.0,0.0078125,-0.0078125,-0.03125,-0.0546875,-0.0234375,-0.0,-0.0234375,0.0078125,-0.0390625,-0.015625,-0.0078125,-0.0390625,0.0234375,-0.0,0.0625,-0.0078125,0.0,0.0390625,0.015625,-0.03125,0.0078125,-0.015625,-0.0078125,0.0625,-0.0546875,-0.03125,0.0234375,0.0625,0.015625,-0.109375,-0.0,-0.0390625,-0.015625,-0.0546875,-0.0078125,-0.0859375,-0.03125,-0.0546875,0.0625,0.0,-0.03125,-0.0078125,-0.0234375,0.0,0.0078125,-0.0078125,-0.0078125,0.03125,0.0078125,-0.0,-0.046875,-0.0546875,0.0,0.0234375,-0.015625,-0.0078125,0.0234375,0.0625,0.0078125,-0.0703125,-0.046875,-0.015625,0.0625,-0.0390625,-0.0234375,-0.0234375,0.0390625,-0.0234375,0.0,0.015625,-0.03125,-0.03125,-0.1015625,-0.03125,-0.0234375,-0.0625,-0.03125,-0.0,-0.109375,-0.0078125,-0.0078125,-0.03125,0.0234375,-0.046875,0.1015625,0.015625,-0.03125,-0.0546875,-0.015625,-0.03125,0.0078125,0.0234375,0.125,-0.0234375,-0.03125,-0.0078125,-0.03125,-0.0390625,0.0625,-0.0390625,0.0234375,0.0234375,-0.0390625,-0.0078125,-0.046875,0.0546875,-0.03125,0.0859375,-0.015625,-0.078125,-0.03125,-0.03125,-0.0234375,-0.0625,-0.0625,-0.015625,0.03125,0.0390625,0.0078125,0.0234375,0.015625,0.0234375,-0.0078125,0.0625,-0.015625,0.0,-0.0546875,0.03125,0.0,0.03125,0.0,0.0234375,-0.0078125,-0.0,-0.0625,-0.0234375,-0.015625,0.0234375,-0.03125,-0.0546875,0.0703125,-0.0078125,-0.046875,0.078125,0.0390625,-0.0625,-0.09375,-0.0546875,0.03125,0.046875,-0.0234375,-0.0078125,-0.0390625,-0.0390625,-0.0078125,0.078125,-0.0078125,0.0234375,-0.0078125,0.0078125,-0.0,-0.0390625,-0.0,-0.0234375,-0.03125,0.0,-0.0234375,-0.03125,0.0546875,-0.0234375,-0.03125,-0.0546875,-0.046875,0.015625,0.0625,-0.03125,-0.03125,0.09375,0.015625,0.046875,-0.0390625,-0.015625,-0.0078125,-0.0625,-0.015625];


outputs = [0.125,0.1875,0.3125,0.125,0.125,0.1875,0.3125,0.125,0.125,0.25,0.125,0.0625,0.1875,0.1875,0.1875,0.0,0.0,0.0,0.0,0.0,0.0,0.0625,0.125,0.0,0.0,0.0,0.0625,0.3125,0.25,0.5,0.3125,0.0625,0.375,0.0625,0.0,0.0625,0.0,0.0,0.0,0.0625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.125,0.0,0.0625,0.4375,0.125,0.125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0625,0.0625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.125,0.0625,0.0,0.0,0.0,0.0,0.0,0.0,0.4375,0.1875,0.25,0.0,0.0,0.0,0.1875,0.0,0.0,0.1875,0.0625,0.125,0.0,0.0,0.25,0.0,0.0,0.0,0.4375,0.0,0.375,0.1875,0.125,0.125,0.3125,0.0625,0.1875,0.375,0.1875,0.25,0.0,0.0,0.0,0.0,0.3125,0.1875,0.0,0.25,0.25,0.25,0.4375,0.5,0.375,0.1875,0.1875,0.1875,0.0,0.0,0.125,0.0625,0.0625,0.0625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.5625,0.125,0.375,0.1875,0.1875,0.25,0.125,0.0625,0.25,0.0,0.0,0.0,0.25,0.0,0.0625,0.125,0.0,0.1875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.125,0.0,0.3125,0.125,0.3125,0.3125,0.0,0.3125,0.5,0.0625,0.3125,0.125,0.125,0.3125,0.0,0.0,0.1875,0.5,0.0625,0.3125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0625,0.0,0.0,0.0,0.0,0.0,0.1875,0.3125,0.0,0.0,0.0,0.0,0.125,0.0,0.375,0.1875,0.25,0.1875,0.0,0.1875,0.0,0.0,0.0,0.125,0.0,0.0625,0.0,0.0625,0.0,0.0,0.0,0.0,0.125,0.1875,0.125,0.125,0.125,0.0625,0.0,0.0625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0625,0.0,0.0,0.0625,0.0,0.4375,0.4375,0.5,0.5,0.0625,0.25,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0625,0.0,0.0,0.125,0.125,0.0625,0.0625,0.0625,0.1875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1875,0.0,0.0625,0.125,0.1875,0.0625,0.0,0.0,0.0,0.0,0.0625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1875,0.1875,0.0625,0.0625,0.0625,0.0,0.0,0.0,0.0,0.375,0.25,0.875,0.125,0.0,0.375,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0625,0.1875,0.25,0.3125,0.3125,0.5,0.125,0.375,0.5,0.0,0.5,0.4375,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.125,0.0,0.0,0.3125,0.375,0.0,0.0,0.1875,0.375,0.0625,0.0625,0.375,0.5,0.375,0.25,0.1875,0.375,0.0,0.0625,0.0625,0.0,0.0,0.1875,0.0,0.0,0.0,0.0,0.0,0.0,0.3125,0.4375,0.1875,0.1875,0.1875,0.375,0.0,0.0,0.0,0.3125,0.125,0.125,0.0625,0.0,0.0,0.125,0.25,0.0,0.4375,0.5,0.5,0.0,0.25,0.4375,0.0,0.0,0.0,0.5625,0.125,0.0,0.0625,0.125,0.125,0.3125,0.375,0.3125,0.375,0.125,0.25,0.1875,0.0,0.0625,0.0,0.0625,0.0,0.1875,0.375,0.125,0.125,0.125,0.1875,0.1875,0.25,0.25,0.0,0.0,0.0,0.0,0.25,0.0,0.1875,0.375,0.3125,0.1875,0.25,0.3125,0.0625,0.0625,0.375,0.3125,0.0,0.1875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.3125,0.125,0.0,0.125,0.0625,0.0625,0.375,0.25,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0625,0.0,0.0,0.0,0.0,0.125,0.0,0.0,0.0,0.1875,0.3125,0.0,0.0,0.1875,0.0,0.0,0.0,0.0,0.125,0.0625,0.0625,0.0,0.0625,0.3125,0.125,0.375,0.0625,0.1875,0.3125,0.0,0.0625,0.0,0.0,0.0,0.375,0.0,0.0,0.0625,0.0,0.0625,0.0,0.0,0.0,0.0,0.0,0.0625,0.0,0.0,0.375,0.1875,0.0625,0.0625,0.0,0.0,0.0,0.0625,0.125,0.0,0.0625,0.0625,0.0,0.1875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.125,0.0,0.0,0.0,0.0,0.0,0.6875,0.125,0.0625,0.4375,0.0,0.0625,0.625,0.0625,0.25,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0625,0.1875,0.0,0.0,0.0,0.0,0.25,0.125,0.125,0.125,0.25,0.0625,0.125,0.1875,0.0,0.0625,0.1875,0.0,0.0,0.0625,0.125,0.0625,0.0,0.0,0.0,0.0,0.3125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0625,0.125,0.0,0.0,0.0625,0.0625,0.0,0.0625,0.3125,0.0625,0.3125,0.6875,0.125,0.5625,0.3125,0.0625,0.3125,0.0,0.0625,0.0,0.125,0.0625,0.25,0.0,0.0,0.0625,0.0,0.0,0.0,0.1875,0.0,0.0,0.0625,0.0625,0.0625,0.4375,0.375,0.4375,0.0,0.0,0.0,0.0625,0.0625,0.0625,0.0,0.0,0.0,0.3125,0.125,0.3125,0.1875,0.0625,0.125,0.125,0.0,0.125,0.5625,0.3125,0.375,0.4375,0.125,0.375,0.4375,0.3125,0.5,0.4375,0.25,0.375,0.3125,0.0,0.1875,0.0,0.0,0.0,0.0,0.0,0.125,0.0,0.0,0.0625,0.0,0.0,0.0,0.0,0.125,0.0,0.0,0.25,0.1875,0.4375,0.1875,0.5,0.4375,0.0,0.625,0.5625,0.0625,0.375,0.6875,0.1875,0.375,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.5625,0.0625,0.1875,0.4375,0.0,0.1875,0.125,0.375,0.375,0.6875,0.0,0.0625,0.25,0.125,0.125,0.125,0.6875,0.4375,0.75,0.5625,0.0,0.5,0.375,0.0625,0.125,0.0,0.0,0.0,0.0,0.0,0.0,0.25,0.3125,0.125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0625,0.1875,0.5625,0.0,0.0,0.0,0.0,0.0,0.0,0.1875,0.0625,0.3125,0.0625,0.0,0.125,0.0,0.0,0.0,0.3125,0.375,0.8125,0.4375,0.0,0.5,0.0,0.0,0.0,0.125,0.0625,0.0,0.0625,0.1875,0.0,0.3125,0.25,0.25,0.125,0.125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0625,0.0,0.0625,0.125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.125,0.0,0.0,0.0,0.25,0.0,0.0,0.0,0.0,0.0,0.0,0.125,0.0,0.0,0.0625,0.1875,0.0,0.125,0.1875,0.25,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.3125,0.4375,0.375,0.25,0.125,0.5625,0.375,0.125,0.4375,0.3125,0.1875,0.0,0.1875,0.125,0.0,0.5,0.0625,0.125,0.8125,0.5625,0.8125,1.25,0.1875,0.6875,0.0625,0.0,0.0,0.125,0.0,0.0,0.125,0.0,0.0,0.125,0.0,0.0,0.0,0.1875,0.375,0.0,0.0,0.25,0.0,0.1875,0.25,0.125,0.0,0.0,0.0625,0.125,0.0625,0.1875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.125,0.0625,0.0,0.0,0.0,0.0,0.0,0.0,0.75,0.125,0.5,0.0,0.0625,0.0625,0.0,0.0,0.0,0.0,0.0,0.0,0.375,0.0,0.25,0.1875,0.0,0.0,0.75,0.375,0.5,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0625,0.0625,0.125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0625,0.0,0.0,0.0,0.0625,0.0,0.1875,0.1875,0.0625,0.0,0.0,0.0,0.0,0.0625,0.0625,0.125,0.25,0.4375,0.1875,0.0625,0.0,0.125,0.0,0.0,0.0,0.0,0.0,0.1875,0.1875,0.5625,0.0,0.0,0.0,0.3125,0.125,0.0,0.0,0.125,0.0,0.0625,0.0,0.0,0.125,0.125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1875,0.125,0.25,0.375,0.125,0.6875,0.375,0.0,0.125,0.3125,0.125,0.0,0.3125,0.0,0.1875,0.125,0.0625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.125,0.0625,0.0,0.0,0.0,0.0,0.0625,0.1875,0.1875,0.125,0.1875,0.125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1875,0.1875,0.1875,0.0,0.0,0.125,0.4375,0.1875,0.5,0.0,0.0,0.0,0.0,0.0625,0.125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.5,0.25,0.375,0.5,0.375,0.75,0.25,0.0625,0.75,0.0,0.0,0.0,0.1875,0.0,0.0,0.4375,0.0,0.0,0.3125,0.0,0.0,0.0,0.0,0.25,0.0,0.0,0.0,0.4375,0.0,0.0,0.375,0.125,0.0625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0625,0.0,0.0,0.1875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.125,0.375,0.0,0.0,0.0,0.375,0.0,0.9375,1.4375,0.1875,0.0,0.3125,0.0,0.0,0.0,0.0,0.0,0.4375,0.875,0.0,0.5,0.5,0.4375,0.25,0.25,0.0,0.625,0.0,0.1875,0.1875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.4375,0.0625,0.375,0.0625,0.0,0.0,0.5625,0.0,0.3125,0.25,0.0,0.125,0.125,0.375,0.5,0.0,0.0,0.3125,0.0625,0.0,0.5,0.0,0.0,0.0,0.5625,0.125,0.125,0.125,0.0625,0.0,0.125,0.0,0.6875,0.0,0.0,0.0,0.5625,0.0,0.1875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.125,0.0,0.0,0.0,0.0,0.0,0.0,0.1875,1.125,0.25,0.0,0.0,0.0625,0.0,0.0,0.0,0.0,0.0,0.1875,0.0,0.3125,0.0,0.3125,1.375,0.0,0.0,0.0,0.0,0.3125,0.0,0.0,0.375,0.0,0.0,0.0,0.0,0.0,0.125,0.0625,0.0,0.0,0.1875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1875,0.25,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.3125,0.0,0.25,0.1875,0.1875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0625,0.0,0.0,0.0625,0.25,0.125,0.3125,0.625,0.0,0.0,0.375,0.0,0.0,0.0,0.0,0.0,0.125,0.25,0.0,0.1875,0.3125,0.1875,0.5,0.4375,0.0,0.75,0.5625,0.0,0.0,0.75,0.125,0.0625,0.0,0.0,0.0,0.0,0.125,0.0,0.0,0.875,0.0,0.0,0.0,0.0,0.0,0.0625,0.0,0.25,0.25,0.0,0.0,0.0,0.0,0.125,0.0,0.125,0.625,0.0,0.3125,1.0,0.0,0.0,0.1875,0.0,0.0,0.0,0.0,0.1875,0.0,0.125,0.75,0.0,0.0,0.0,0.375,0.0625,0.5,0.375,0.0,0.1875,0.0,0.0,0.0625,0.0,0.0,0.0,0.0,0.0,0.375,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.375,0.125,0.0,0.0,0.0,0.0,0.0,0.0,0.5625,0.0,0.0,0.375,0.0,0.0625,0.0,0.0,0.0,0.0,0.5,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0625,0.0,0.0,0.1875,0.0,0.0625,0.3125,0.0,0.0,0.0,0.0,0.0,0.0,0.6875,0.0,0.0,0.0,0.0,0.3125,0.9375,1.5,0.0,0.0,0.1875,0.6875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.125,0.0,0.1875,0.0625,0.0,0.0,0.0,0.0,0.0,0.6875,0.3125,0.0,0.0,0.0,0.0,0.5,0.875,0.4375,0.3125,0.5,0.0,0.0,0.1875,0.6875,0.125,0.6875,0.0,0.25,0.5625,0.6875,0.1875,0.625,0.125,0.0,0.1875,0.0,0.125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.125,0.0,0.0,0.75,0.0,0.0,0.0,0.0,0.0,0.0625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.3125,0.0,0.0,0.0625,0.0,0.0,0.0,0.0,0.0,0.25,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.25,0.1875,0.0,0.375,0.8125,0.4375,0.0,0.25,0.0625,0.0,0.0,0.0,0.0,0.0,0.0,0.1875,0.0,0.25,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.125,0.125,0.0,0.5625,0.0625,0.0,0.0,0.0,0.0,0.0,0.375,0.0625,0.5,0.0,0.1875,0.0,0.0,0.0,0.0,0.4375,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.875,0.0,0.0,0.0,0.375,0.0,0.0,0.1875,0.0625,0.0625,0.0625,0.125,0.25,0.75,0.25,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.4375,0.6875,0.625,0.6875,0.75,0.0,0.0,0.0,0.0,0.0,0.0,0.1875,0.0,0.0,0.375,0.75,0.1875,0.0,0.1875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.125,0.0,0.0,0.125,0.0,0.0,0.0625,0.0625,0.9375,0.0,0.0,0.8125,0.0,0.0,0.4375,0.0,0.0625,0.0,0.0,0.8125,0.0,0.0,0.3125,0.25,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.25,0.25,0.0,0.0,0.0,0.0,0.5625,0.0,0.5,0.75,0.0,0.5625,0.0,0.0,0.0,0.0,0.0625,0.0,0.0,0.0,0.0,0.6875,0.0,0.0,0.1875,0.0,0.0,0.0,0.375,0.0,0.1875,0.4375,0.25,0.0,0.0,0.0,0.0,0.25,0.0,0.25,1.0625,0.1875,0.75,1.4375,0.5,0.0,0.0,0.0,0.0,0.1875,0.0625,0.0,0.0,0.0,0.1875,0.125,0.125,0.0,0.0,0.0,0.0,0.0,0.0625,0.0,0.0,0.0,0.125,0.0,0.0,0.0,0.0,0.125,0.0,0.0,0.0625,0.0,0.0,0.0,0.0,0.0,0.0,0.375,0.0,0.0,0.3125,1.3125,0.375,0.0,1.0,0.0,0.0,0.6875,0.0,0.0,0.0,0.0,0.0625,0.0,0.0,0.1875,0.0,0.125,0.0,0.0,0.0,0.0,0.0,0.0,0.0625,0.3125,0.0,0.125,0.0,0.0,0.5,0.8125,0.9375,0.8125,0.1875,0.8125,0.5,0.5,0.8125,0.0,0.0,0.0,0.8125,0.0,0.4375,0.0,0.0,0.0,0.0,0.0,0.125,0.0,0.5625,0.6875,0.0,0.3125,0.0,0.0,0.0,0.125,0.0,0.0625,0.3125,0.25,0.4375,0.5,0.0,0.0,0.0,0.1875,0.0,0.25,0.0,0.0,0.0,0.1875,0.1875,0.0,0.0,0.4375,0.0,0.375,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.75,0.0,0.4375,0.3125,0.0,0.125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.0,0.3125,0.75,0.9375,0.0,1.1875,1.1875,1.125,0.9375,0.0,0.0,0.0,0.0,1.4375,1.0625,0.0,0.0625,0.5,0.1875,0.125,0.0,0.0625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.5,0.625,0.25,1.0,0.5625,0.0,0.0625,0.25,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.5625,0.3125,0.0,0.0,0.1875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.375,0.0,0.0625,0.25,0.4375,0.8125,0.9375,0.75,0.5625,0.125,0.375,0.0,0.0,0.0,0.0,0.8125,0.0,0.0,1.0625,0.0,0.0,0.9375,0.0,0.0,0.0,0.0625,0.0,0.0,0.1875,0.25,0.0,0.0,0.25,0.0,0.0,0.0,0.0,0.0,0.0,0.0625,0.0,0.4375,0.0,0.5,0.5625,0.0,0.8125,0.3125,0.125,0.25,0.0,0.0,0.0,0.0,0.9375,0.0,0.0,0.0,0.0,0.6875,0.0,0.6875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.25,0.0,0.375,0.75,0.0,0.4375,0.0,0.75,0.0,0.4375,0.875,0.5625,0.0,0.0,0.0625,0.0,0.0625,0.75,0.0,0.0,0.0,0.0625,0.1875,0.0,0.0,0.0,0.0,0.75,1.125,0.6875,0.0,0.0,0.0,0.125,0.3125,0.0,0.0625,0.0625,0.0,0.0625,0.0,0.125,0.0,0.0,0.0,0.4375,0.0,0.3125,0.0,0.0,0.0,0.4375,0.3125,1.0625,0.0,0.0,0.8125,0.5,0.0625,0.75,0.25,0.5,0.3125,0.0,0.0,0.0,0.125,0.0,0.25,0.1875,0.0,0.0,0.5625,0.0,0.0,0.0,0.8125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1875,0.0,0.0,0.4375,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.25,0.0,0.0,0.125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.5,0.25,0.4375,0.0,0.5625,0.625,0.375,1.3125,0.125,0.5625,0.6875,0.25,0.0,0.0,0.0,0.375,0.0625,0.125,0.375,0.1875,0.5625,0.0,0.0,0.0,0.5,0.0,0.8125,0.5,0.0625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.4375,0.3125,0.0625,0.625];



endpackage : arrays